library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package TXT_LIB is

	type CoordPair is record
	  x : integer; 
	  y : integer;
	end record;
	type CoordPairArray is array (natural range <>) of CoordPair;
	
	constant start_screen_arr: CoordPairArray(0 to 4449) := (
  (x => 293, y => 151),
  (x => 294, y => 151),
  (x => 295, y => 151),
  (x => 296, y => 151),
  (x => 297, y => 151),
  (x => 298, y => 151),
  (x => 299, y => 151),
  (x => 300, y => 151),
  (x => 301, y => 151),
  (x => 302, y => 151),
  (x => 379, y => 151),
  (x => 380, y => 151),
  (x => 381, y => 151),
  (x => 382, y => 151),
  (x => 383, y => 151),
  (x => 384, y => 151),
  (x => 385, y => 151),
  (x => 386, y => 151),
  (x => 387, y => 151),
  (x => 388, y => 151),
  (x => 389, y => 151),
  (x => 249, y => 152),
  (x => 250, y => 152),
  (x => 251, y => 152),
  (x => 252, y => 152),
  (x => 253, y => 152),
  (x => 254, y => 152),
  (x => 255, y => 152),
  (x => 256, y => 152),
  (x => 257, y => 152),
  (x => 258, y => 152),
  (x => 259, y => 152),
  (x => 260, y => 152),
  (x => 261, y => 152),
  (x => 262, y => 152),
  (x => 263, y => 152),
  (x => 264, y => 152),
  (x => 265, y => 152),
  (x => 266, y => 152),
  (x => 291, y => 152),
  (x => 292, y => 152),
  (x => 293, y => 152),
  (x => 294, y => 152),
  (x => 295, y => 152),
  (x => 296, y => 152),
  (x => 297, y => 152),
  (x => 298, y => 152),
  (x => 299, y => 152),
  (x => 300, y => 152),
  (x => 301, y => 152),
  (x => 302, y => 152),
  (x => 303, y => 152),
  (x => 304, y => 152),
  (x => 323, y => 152),
  (x => 324, y => 152),
  (x => 325, y => 152),
  (x => 326, y => 152),
  (x => 327, y => 152),
  (x => 328, y => 152),
  (x => 329, y => 152),
  (x => 330, y => 152),
  (x => 331, y => 152),
  (x => 349, y => 152),
  (x => 350, y => 152),
  (x => 351, y => 152),
  (x => 352, y => 152),
  (x => 353, y => 152),
  (x => 354, y => 152),
  (x => 355, y => 152),
  (x => 376, y => 152),
  (x => 377, y => 152),
  (x => 378, y => 152),
  (x => 379, y => 152),
  (x => 380, y => 152),
  (x => 381, y => 152),
  (x => 382, y => 152),
  (x => 383, y => 152),
  (x => 384, y => 152),
  (x => 385, y => 152),
  (x => 386, y => 152),
  (x => 387, y => 152),
  (x => 388, y => 152),
  (x => 389, y => 152),
  (x => 390, y => 152),
  (x => 391, y => 152),
  (x => 392, y => 152),
  (x => 249, y => 153),
  (x => 250, y => 153),
  (x => 251, y => 153),
  (x => 252, y => 153),
  (x => 253, y => 153),
  (x => 254, y => 153),
  (x => 255, y => 153),
  (x => 256, y => 153),
  (x => 257, y => 153),
  (x => 258, y => 153),
  (x => 259, y => 153),
  (x => 260, y => 153),
  (x => 261, y => 153),
  (x => 262, y => 153),
  (x => 263, y => 153),
  (x => 264, y => 153),
  (x => 265, y => 153),
  (x => 266, y => 153),
  (x => 267, y => 153),
  (x => 268, y => 153),
  (x => 269, y => 153),
  (x => 289, y => 153),
  (x => 290, y => 153),
  (x => 291, y => 153),
  (x => 292, y => 153),
  (x => 293, y => 153),
  (x => 294, y => 153),
  (x => 295, y => 153),
  (x => 296, y => 153),
  (x => 297, y => 153),
  (x => 298, y => 153),
  (x => 299, y => 153),
  (x => 300, y => 153),
  (x => 301, y => 153),
  (x => 302, y => 153),
  (x => 303, y => 153),
  (x => 304, y => 153),
  (x => 305, y => 153),
  (x => 306, y => 153),
  (x => 323, y => 153),
  (x => 324, y => 153),
  (x => 325, y => 153),
  (x => 326, y => 153),
  (x => 327, y => 153),
  (x => 328, y => 153),
  (x => 329, y => 153),
  (x => 330, y => 153),
  (x => 331, y => 153),
  (x => 349, y => 153),
  (x => 350, y => 153),
  (x => 351, y => 153),
  (x => 352, y => 153),
  (x => 353, y => 153),
  (x => 354, y => 153),
  (x => 355, y => 153),
  (x => 374, y => 153),
  (x => 375, y => 153),
  (x => 376, y => 153),
  (x => 377, y => 153),
  (x => 378, y => 153),
  (x => 379, y => 153),
  (x => 380, y => 153),
  (x => 381, y => 153),
  (x => 382, y => 153),
  (x => 383, y => 153),
  (x => 384, y => 153),
  (x => 385, y => 153),
  (x => 386, y => 153),
  (x => 387, y => 153),
  (x => 388, y => 153),
  (x => 389, y => 153),
  (x => 390, y => 153),
  (x => 391, y => 153),
  (x => 392, y => 153),
  (x => 393, y => 153),
  (x => 249, y => 154),
  (x => 250, y => 154),
  (x => 251, y => 154),
  (x => 252, y => 154),
  (x => 253, y => 154),
  (x => 254, y => 154),
  (x => 255, y => 154),
  (x => 256, y => 154),
  (x => 257, y => 154),
  (x => 258, y => 154),
  (x => 259, y => 154),
  (x => 260, y => 154),
  (x => 261, y => 154),
  (x => 262, y => 154),
  (x => 263, y => 154),
  (x => 264, y => 154),
  (x => 265, y => 154),
  (x => 266, y => 154),
  (x => 267, y => 154),
  (x => 268, y => 154),
  (x => 269, y => 154),
  (x => 270, y => 154),
  (x => 288, y => 154),
  (x => 289, y => 154),
  (x => 290, y => 154),
  (x => 291, y => 154),
  (x => 292, y => 154),
  (x => 293, y => 154),
  (x => 294, y => 154),
  (x => 295, y => 154),
  (x => 296, y => 154),
  (x => 297, y => 154),
  (x => 298, y => 154),
  (x => 299, y => 154),
  (x => 300, y => 154),
  (x => 301, y => 154),
  (x => 302, y => 154),
  (x => 303, y => 154),
  (x => 304, y => 154),
  (x => 305, y => 154),
  (x => 306, y => 154),
  (x => 307, y => 154),
  (x => 323, y => 154),
  (x => 324, y => 154),
  (x => 325, y => 154),
  (x => 326, y => 154),
  (x => 327, y => 154),
  (x => 328, y => 154),
  (x => 329, y => 154),
  (x => 330, y => 154),
  (x => 331, y => 154),
  (x => 332, y => 154),
  (x => 349, y => 154),
  (x => 350, y => 154),
  (x => 351, y => 154),
  (x => 352, y => 154),
  (x => 353, y => 154),
  (x => 354, y => 154),
  (x => 355, y => 154),
  (x => 373, y => 154),
  (x => 374, y => 154),
  (x => 375, y => 154),
  (x => 376, y => 154),
  (x => 377, y => 154),
  (x => 378, y => 154),
  (x => 379, y => 154),
  (x => 380, y => 154),
  (x => 381, y => 154),
  (x => 382, y => 154),
  (x => 383, y => 154),
  (x => 384, y => 154),
  (x => 385, y => 154),
  (x => 386, y => 154),
  (x => 387, y => 154),
  (x => 388, y => 154),
  (x => 389, y => 154),
  (x => 390, y => 154),
  (x => 391, y => 154),
  (x => 392, y => 154),
  (x => 393, y => 154),
  (x => 249, y => 155),
  (x => 250, y => 155),
  (x => 251, y => 155),
  (x => 252, y => 155),
  (x => 253, y => 155),
  (x => 254, y => 155),
  (x => 255, y => 155),
  (x => 256, y => 155),
  (x => 257, y => 155),
  (x => 258, y => 155),
  (x => 259, y => 155),
  (x => 260, y => 155),
  (x => 261, y => 155),
  (x => 262, y => 155),
  (x => 263, y => 155),
  (x => 264, y => 155),
  (x => 265, y => 155),
  (x => 266, y => 155),
  (x => 267, y => 155),
  (x => 268, y => 155),
  (x => 269, y => 155),
  (x => 270, y => 155),
  (x => 271, y => 155),
  (x => 287, y => 155),
  (x => 288, y => 155),
  (x => 289, y => 155),
  (x => 290, y => 155),
  (x => 291, y => 155),
  (x => 292, y => 155),
  (x => 293, y => 155),
  (x => 294, y => 155),
  (x => 295, y => 155),
  (x => 296, y => 155),
  (x => 297, y => 155),
  (x => 298, y => 155),
  (x => 299, y => 155),
  (x => 300, y => 155),
  (x => 301, y => 155),
  (x => 302, y => 155),
  (x => 303, y => 155),
  (x => 304, y => 155),
  (x => 305, y => 155),
  (x => 306, y => 155),
  (x => 307, y => 155),
  (x => 308, y => 155),
  (x => 323, y => 155),
  (x => 324, y => 155),
  (x => 325, y => 155),
  (x => 326, y => 155),
  (x => 327, y => 155),
  (x => 328, y => 155),
  (x => 329, y => 155),
  (x => 330, y => 155),
  (x => 331, y => 155),
  (x => 332, y => 155),
  (x => 349, y => 155),
  (x => 350, y => 155),
  (x => 351, y => 155),
  (x => 352, y => 155),
  (x => 353, y => 155),
  (x => 354, y => 155),
  (x => 355, y => 155),
  (x => 371, y => 155),
  (x => 372, y => 155),
  (x => 373, y => 155),
  (x => 374, y => 155),
  (x => 375, y => 155),
  (x => 376, y => 155),
  (x => 377, y => 155),
  (x => 378, y => 155),
  (x => 379, y => 155),
  (x => 380, y => 155),
  (x => 381, y => 155),
  (x => 382, y => 155),
  (x => 383, y => 155),
  (x => 384, y => 155),
  (x => 385, y => 155),
  (x => 386, y => 155),
  (x => 387, y => 155),
  (x => 388, y => 155),
  (x => 389, y => 155),
  (x => 390, y => 155),
  (x => 391, y => 155),
  (x => 392, y => 155),
  (x => 393, y => 155),
  (x => 249, y => 156),
  (x => 250, y => 156),
  (x => 251, y => 156),
  (x => 252, y => 156),
  (x => 253, y => 156),
  (x => 254, y => 156),
  (x => 255, y => 156),
  (x => 256, y => 156),
  (x => 257, y => 156),
  (x => 258, y => 156),
  (x => 259, y => 156),
  (x => 260, y => 156),
  (x => 261, y => 156),
  (x => 262, y => 156),
  (x => 263, y => 156),
  (x => 264, y => 156),
  (x => 265, y => 156),
  (x => 266, y => 156),
  (x => 267, y => 156),
  (x => 268, y => 156),
  (x => 269, y => 156),
  (x => 270, y => 156),
  (x => 271, y => 156),
  (x => 272, y => 156),
  (x => 286, y => 156),
  (x => 287, y => 156),
  (x => 288, y => 156),
  (x => 289, y => 156),
  (x => 290, y => 156),
  (x => 291, y => 156),
  (x => 292, y => 156),
  (x => 293, y => 156),
  (x => 294, y => 156),
  (x => 295, y => 156),
  (x => 296, y => 156),
  (x => 297, y => 156),
  (x => 298, y => 156),
  (x => 299, y => 156),
  (x => 300, y => 156),
  (x => 301, y => 156),
  (x => 302, y => 156),
  (x => 303, y => 156),
  (x => 304, y => 156),
  (x => 305, y => 156),
  (x => 306, y => 156),
  (x => 307, y => 156),
  (x => 308, y => 156),
  (x => 309, y => 156),
  (x => 323, y => 156),
  (x => 324, y => 156),
  (x => 325, y => 156),
  (x => 326, y => 156),
  (x => 327, y => 156),
  (x => 328, y => 156),
  (x => 329, y => 156),
  (x => 330, y => 156),
  (x => 331, y => 156),
  (x => 332, y => 156),
  (x => 333, y => 156),
  (x => 349, y => 156),
  (x => 350, y => 156),
  (x => 351, y => 156),
  (x => 352, y => 156),
  (x => 353, y => 156),
  (x => 354, y => 156),
  (x => 355, y => 156),
  (x => 371, y => 156),
  (x => 372, y => 156),
  (x => 373, y => 156),
  (x => 374, y => 156),
  (x => 375, y => 156),
  (x => 376, y => 156),
  (x => 377, y => 156),
  (x => 378, y => 156),
  (x => 379, y => 156),
  (x => 380, y => 156),
  (x => 381, y => 156),
  (x => 382, y => 156),
  (x => 383, y => 156),
  (x => 384, y => 156),
  (x => 385, y => 156),
  (x => 386, y => 156),
  (x => 387, y => 156),
  (x => 388, y => 156),
  (x => 389, y => 156),
  (x => 390, y => 156),
  (x => 391, y => 156),
  (x => 392, y => 156),
  (x => 393, y => 156),
  (x => 249, y => 157),
  (x => 250, y => 157),
  (x => 251, y => 157),
  (x => 252, y => 157),
  (x => 253, y => 157),
  (x => 254, y => 157),
  (x => 255, y => 157),
  (x => 256, y => 157),
  (x => 257, y => 157),
  (x => 258, y => 157),
  (x => 259, y => 157),
  (x => 260, y => 157),
  (x => 261, y => 157),
  (x => 262, y => 157),
  (x => 263, y => 157),
  (x => 264, y => 157),
  (x => 265, y => 157),
  (x => 266, y => 157),
  (x => 267, y => 157),
  (x => 268, y => 157),
  (x => 269, y => 157),
  (x => 270, y => 157),
  (x => 271, y => 157),
  (x => 272, y => 157),
  (x => 273, y => 157),
  (x => 285, y => 157),
  (x => 286, y => 157),
  (x => 287, y => 157),
  (x => 288, y => 157),
  (x => 289, y => 157),
  (x => 290, y => 157),
  (x => 291, y => 157),
  (x => 292, y => 157),
  (x => 293, y => 157),
  (x => 294, y => 157),
  (x => 295, y => 157),
  (x => 296, y => 157),
  (x => 297, y => 157),
  (x => 298, y => 157),
  (x => 299, y => 157),
  (x => 300, y => 157),
  (x => 301, y => 157),
  (x => 302, y => 157),
  (x => 303, y => 157),
  (x => 304, y => 157),
  (x => 305, y => 157),
  (x => 306, y => 157),
  (x => 307, y => 157),
  (x => 308, y => 157),
  (x => 309, y => 157),
  (x => 310, y => 157),
  (x => 323, y => 157),
  (x => 324, y => 157),
  (x => 325, y => 157),
  (x => 326, y => 157),
  (x => 327, y => 157),
  (x => 328, y => 157),
  (x => 329, y => 157),
  (x => 330, y => 157),
  (x => 331, y => 157),
  (x => 332, y => 157),
  (x => 333, y => 157),
  (x => 349, y => 157),
  (x => 350, y => 157),
  (x => 351, y => 157),
  (x => 352, y => 157),
  (x => 353, y => 157),
  (x => 354, y => 157),
  (x => 355, y => 157),
  (x => 370, y => 157),
  (x => 371, y => 157),
  (x => 372, y => 157),
  (x => 373, y => 157),
  (x => 374, y => 157),
  (x => 375, y => 157),
  (x => 376, y => 157),
  (x => 377, y => 157),
  (x => 378, y => 157),
  (x => 379, y => 157),
  (x => 380, y => 157),
  (x => 381, y => 157),
  (x => 382, y => 157),
  (x => 383, y => 157),
  (x => 384, y => 157),
  (x => 385, y => 157),
  (x => 386, y => 157),
  (x => 387, y => 157),
  (x => 388, y => 157),
  (x => 389, y => 157),
  (x => 390, y => 157),
  (x => 391, y => 157),
  (x => 392, y => 157),
  (x => 393, y => 157),
  (x => 249, y => 158),
  (x => 250, y => 158),
  (x => 251, y => 158),
  (x => 252, y => 158),
  (x => 253, y => 158),
  (x => 254, y => 158),
  (x => 255, y => 158),
  (x => 256, y => 158),
  (x => 257, y => 158),
  (x => 258, y => 158),
  (x => 259, y => 158),
  (x => 260, y => 158),
  (x => 261, y => 158),
  (x => 262, y => 158),
  (x => 263, y => 158),
  (x => 264, y => 158),
  (x => 265, y => 158),
  (x => 266, y => 158),
  (x => 267, y => 158),
  (x => 268, y => 158),
  (x => 269, y => 158),
  (x => 270, y => 158),
  (x => 271, y => 158),
  (x => 272, y => 158),
  (x => 273, y => 158),
  (x => 285, y => 158),
  (x => 286, y => 158),
  (x => 287, y => 158),
  (x => 288, y => 158),
  (x => 289, y => 158),
  (x => 290, y => 158),
  (x => 291, y => 158),
  (x => 292, y => 158),
  (x => 293, y => 158),
  (x => 294, y => 158),
  (x => 295, y => 158),
  (x => 296, y => 158),
  (x => 297, y => 158),
  (x => 298, y => 158),
  (x => 299, y => 158),
  (x => 300, y => 158),
  (x => 301, y => 158),
  (x => 302, y => 158),
  (x => 303, y => 158),
  (x => 304, y => 158),
  (x => 305, y => 158),
  (x => 306, y => 158),
  (x => 307, y => 158),
  (x => 308, y => 158),
  (x => 309, y => 158),
  (x => 310, y => 158),
  (x => 323, y => 158),
  (x => 324, y => 158),
  (x => 325, y => 158),
  (x => 326, y => 158),
  (x => 327, y => 158),
  (x => 328, y => 158),
  (x => 329, y => 158),
  (x => 330, y => 158),
  (x => 331, y => 158),
  (x => 332, y => 158),
  (x => 333, y => 158),
  (x => 334, y => 158),
  (x => 349, y => 158),
  (x => 350, y => 158),
  (x => 351, y => 158),
  (x => 352, y => 158),
  (x => 353, y => 158),
  (x => 354, y => 158),
  (x => 355, y => 158),
  (x => 369, y => 158),
  (x => 370, y => 158),
  (x => 371, y => 158),
  (x => 372, y => 158),
  (x => 373, y => 158),
  (x => 374, y => 158),
  (x => 375, y => 158),
  (x => 376, y => 158),
  (x => 377, y => 158),
  (x => 378, y => 158),
  (x => 379, y => 158),
  (x => 380, y => 158),
  (x => 381, y => 158),
  (x => 382, y => 158),
  (x => 383, y => 158),
  (x => 384, y => 158),
  (x => 385, y => 158),
  (x => 386, y => 158),
  (x => 387, y => 158),
  (x => 388, y => 158),
  (x => 389, y => 158),
  (x => 390, y => 158),
  (x => 391, y => 158),
  (x => 392, y => 158),
  (x => 393, y => 158),
  (x => 249, y => 159),
  (x => 250, y => 159),
  (x => 251, y => 159),
  (x => 252, y => 159),
  (x => 253, y => 159),
  (x => 254, y => 159),
  (x => 255, y => 159),
  (x => 256, y => 159),
  (x => 264, y => 159),
  (x => 265, y => 159),
  (x => 266, y => 159),
  (x => 267, y => 159),
  (x => 268, y => 159),
  (x => 269, y => 159),
  (x => 270, y => 159),
  (x => 271, y => 159),
  (x => 272, y => 159),
  (x => 273, y => 159),
  (x => 284, y => 159),
  (x => 285, y => 159),
  (x => 286, y => 159),
  (x => 287, y => 159),
  (x => 288, y => 159),
  (x => 289, y => 159),
  (x => 290, y => 159),
  (x => 291, y => 159),
  (x => 292, y => 159),
  (x => 293, y => 159),
  (x => 294, y => 159),
  (x => 301, y => 159),
  (x => 302, y => 159),
  (x => 303, y => 159),
  (x => 304, y => 159),
  (x => 305, y => 159),
  (x => 306, y => 159),
  (x => 307, y => 159),
  (x => 308, y => 159),
  (x => 309, y => 159),
  (x => 310, y => 159),
  (x => 311, y => 159),
  (x => 323, y => 159),
  (x => 324, y => 159),
  (x => 325, y => 159),
  (x => 326, y => 159),
  (x => 327, y => 159),
  (x => 328, y => 159),
  (x => 329, y => 159),
  (x => 330, y => 159),
  (x => 331, y => 159),
  (x => 332, y => 159),
  (x => 333, y => 159),
  (x => 334, y => 159),
  (x => 349, y => 159),
  (x => 350, y => 159),
  (x => 351, y => 159),
  (x => 352, y => 159),
  (x => 353, y => 159),
  (x => 354, y => 159),
  (x => 355, y => 159),
  (x => 368, y => 159),
  (x => 369, y => 159),
  (x => 370, y => 159),
  (x => 371, y => 159),
  (x => 372, y => 159),
  (x => 373, y => 159),
  (x => 374, y => 159),
  (x => 375, y => 159),
  (x => 376, y => 159),
  (x => 377, y => 159),
  (x => 378, y => 159),
  (x => 379, y => 159),
  (x => 390, y => 159),
  (x => 391, y => 159),
  (x => 392, y => 159),
  (x => 393, y => 159),
  (x => 249, y => 160),
  (x => 250, y => 160),
  (x => 251, y => 160),
  (x => 252, y => 160),
  (x => 253, y => 160),
  (x => 254, y => 160),
  (x => 255, y => 160),
  (x => 265, y => 160),
  (x => 266, y => 160),
  (x => 267, y => 160),
  (x => 268, y => 160),
  (x => 269, y => 160),
  (x => 270, y => 160),
  (x => 271, y => 160),
  (x => 272, y => 160),
  (x => 273, y => 160),
  (x => 274, y => 160),
  (x => 284, y => 160),
  (x => 285, y => 160),
  (x => 286, y => 160),
  (x => 287, y => 160),
  (x => 288, y => 160),
  (x => 289, y => 160),
  (x => 290, y => 160),
  (x => 291, y => 160),
  (x => 292, y => 160),
  (x => 303, y => 160),
  (x => 304, y => 160),
  (x => 305, y => 160),
  (x => 306, y => 160),
  (x => 307, y => 160),
  (x => 308, y => 160),
  (x => 309, y => 160),
  (x => 310, y => 160),
  (x => 311, y => 160),
  (x => 312, y => 160),
  (x => 323, y => 160),
  (x => 324, y => 160),
  (x => 325, y => 160),
  (x => 326, y => 160),
  (x => 327, y => 160),
  (x => 328, y => 160),
  (x => 329, y => 160),
  (x => 330, y => 160),
  (x => 331, y => 160),
  (x => 332, y => 160),
  (x => 333, y => 160),
  (x => 334, y => 160),
  (x => 335, y => 160),
  (x => 349, y => 160),
  (x => 350, y => 160),
  (x => 351, y => 160),
  (x => 352, y => 160),
  (x => 353, y => 160),
  (x => 354, y => 160),
  (x => 355, y => 160),
  (x => 368, y => 160),
  (x => 369, y => 160),
  (x => 370, y => 160),
  (x => 371, y => 160),
  (x => 372, y => 160),
  (x => 373, y => 160),
  (x => 374, y => 160),
  (x => 375, y => 160),
  (x => 376, y => 160),
  (x => 377, y => 160),
  (x => 392, y => 160),
  (x => 393, y => 160),
  (x => 249, y => 161),
  (x => 250, y => 161),
  (x => 251, y => 161),
  (x => 252, y => 161),
  (x => 253, y => 161),
  (x => 254, y => 161),
  (x => 255, y => 161),
  (x => 266, y => 161),
  (x => 267, y => 161),
  (x => 268, y => 161),
  (x => 269, y => 161),
  (x => 270, y => 161),
  (x => 271, y => 161),
  (x => 272, y => 161),
  (x => 273, y => 161),
  (x => 274, y => 161),
  (x => 283, y => 161),
  (x => 284, y => 161),
  (x => 285, y => 161),
  (x => 286, y => 161),
  (x => 287, y => 161),
  (x => 288, y => 161),
  (x => 289, y => 161),
  (x => 290, y => 161),
  (x => 291, y => 161),
  (x => 304, y => 161),
  (x => 305, y => 161),
  (x => 306, y => 161),
  (x => 307, y => 161),
  (x => 308, y => 161),
  (x => 309, y => 161),
  (x => 310, y => 161),
  (x => 311, y => 161),
  (x => 312, y => 161),
  (x => 323, y => 161),
  (x => 324, y => 161),
  (x => 325, y => 161),
  (x => 326, y => 161),
  (x => 327, y => 161),
  (x => 328, y => 161),
  (x => 329, y => 161),
  (x => 330, y => 161),
  (x => 331, y => 161),
  (x => 332, y => 161),
  (x => 333, y => 161),
  (x => 334, y => 161),
  (x => 335, y => 161),
  (x => 349, y => 161),
  (x => 350, y => 161),
  (x => 351, y => 161),
  (x => 352, y => 161),
  (x => 353, y => 161),
  (x => 354, y => 161),
  (x => 355, y => 161),
  (x => 367, y => 161),
  (x => 368, y => 161),
  (x => 369, y => 161),
  (x => 370, y => 161),
  (x => 371, y => 161),
  (x => 372, y => 161),
  (x => 373, y => 161),
  (x => 374, y => 161),
  (x => 375, y => 161),
  (x => 376, y => 161),
  (x => 249, y => 162),
  (x => 250, y => 162),
  (x => 251, y => 162),
  (x => 252, y => 162),
  (x => 253, y => 162),
  (x => 254, y => 162),
  (x => 255, y => 162),
  (x => 267, y => 162),
  (x => 268, y => 162),
  (x => 269, y => 162),
  (x => 270, y => 162),
  (x => 271, y => 162),
  (x => 272, y => 162),
  (x => 273, y => 162),
  (x => 274, y => 162),
  (x => 283, y => 162),
  (x => 284, y => 162),
  (x => 285, y => 162),
  (x => 286, y => 162),
  (x => 287, y => 162),
  (x => 288, y => 162),
  (x => 289, y => 162),
  (x => 290, y => 162),
  (x => 305, y => 162),
  (x => 306, y => 162),
  (x => 307, y => 162),
  (x => 308, y => 162),
  (x => 309, y => 162),
  (x => 310, y => 162),
  (x => 311, y => 162),
  (x => 312, y => 162),
  (x => 323, y => 162),
  (x => 324, y => 162),
  (x => 325, y => 162),
  (x => 326, y => 162),
  (x => 327, y => 162),
  (x => 328, y => 162),
  (x => 329, y => 162),
  (x => 330, y => 162),
  (x => 331, y => 162),
  (x => 332, y => 162),
  (x => 333, y => 162),
  (x => 334, y => 162),
  (x => 335, y => 162),
  (x => 336, y => 162),
  (x => 349, y => 162),
  (x => 350, y => 162),
  (x => 351, y => 162),
  (x => 352, y => 162),
  (x => 353, y => 162),
  (x => 354, y => 162),
  (x => 355, y => 162),
  (x => 367, y => 162),
  (x => 368, y => 162),
  (x => 369, y => 162),
  (x => 370, y => 162),
  (x => 371, y => 162),
  (x => 372, y => 162),
  (x => 373, y => 162),
  (x => 374, y => 162),
  (x => 375, y => 162),
  (x => 249, y => 163),
  (x => 250, y => 163),
  (x => 251, y => 163),
  (x => 252, y => 163),
  (x => 253, y => 163),
  (x => 254, y => 163),
  (x => 255, y => 163),
  (x => 267, y => 163),
  (x => 268, y => 163),
  (x => 269, y => 163),
  (x => 270, y => 163),
  (x => 271, y => 163),
  (x => 272, y => 163),
  (x => 273, y => 163),
  (x => 274, y => 163),
  (x => 282, y => 163),
  (x => 283, y => 163),
  (x => 284, y => 163),
  (x => 285, y => 163),
  (x => 286, y => 163),
  (x => 287, y => 163),
  (x => 288, y => 163),
  (x => 289, y => 163),
  (x => 290, y => 163),
  (x => 305, y => 163),
  (x => 306, y => 163),
  (x => 307, y => 163),
  (x => 308, y => 163),
  (x => 309, y => 163),
  (x => 310, y => 163),
  (x => 311, y => 163),
  (x => 312, y => 163),
  (x => 313, y => 163),
  (x => 323, y => 163),
  (x => 324, y => 163),
  (x => 325, y => 163),
  (x => 326, y => 163),
  (x => 327, y => 163),
  (x => 328, y => 163),
  (x => 329, y => 163),
  (x => 330, y => 163),
  (x => 331, y => 163),
  (x => 332, y => 163),
  (x => 333, y => 163),
  (x => 334, y => 163),
  (x => 335, y => 163),
  (x => 336, y => 163),
  (x => 349, y => 163),
  (x => 350, y => 163),
  (x => 351, y => 163),
  (x => 352, y => 163),
  (x => 353, y => 163),
  (x => 354, y => 163),
  (x => 355, y => 163),
  (x => 366, y => 163),
  (x => 367, y => 163),
  (x => 368, y => 163),
  (x => 369, y => 163),
  (x => 370, y => 163),
  (x => 371, y => 163),
  (x => 372, y => 163),
  (x => 373, y => 163),
  (x => 374, y => 163),
  (x => 249, y => 164),
  (x => 250, y => 164),
  (x => 251, y => 164),
  (x => 252, y => 164),
  (x => 253, y => 164),
  (x => 254, y => 164),
  (x => 255, y => 164),
  (x => 268, y => 164),
  (x => 269, y => 164),
  (x => 270, y => 164),
  (x => 271, y => 164),
  (x => 272, y => 164),
  (x => 273, y => 164),
  (x => 274, y => 164),
  (x => 282, y => 164),
  (x => 283, y => 164),
  (x => 284, y => 164),
  (x => 285, y => 164),
  (x => 286, y => 164),
  (x => 287, y => 164),
  (x => 288, y => 164),
  (x => 289, y => 164),
  (x => 306, y => 164),
  (x => 307, y => 164),
  (x => 308, y => 164),
  (x => 309, y => 164),
  (x => 310, y => 164),
  (x => 311, y => 164),
  (x => 312, y => 164),
  (x => 313, y => 164),
  (x => 323, y => 164),
  (x => 324, y => 164),
  (x => 325, y => 164),
  (x => 326, y => 164),
  (x => 327, y => 164),
  (x => 328, y => 164),
  (x => 329, y => 164),
  (x => 330, y => 164),
  (x => 331, y => 164),
  (x => 332, y => 164),
  (x => 333, y => 164),
  (x => 334, y => 164),
  (x => 335, y => 164),
  (x => 336, y => 164),
  (x => 337, y => 164),
  (x => 349, y => 164),
  (x => 350, y => 164),
  (x => 351, y => 164),
  (x => 352, y => 164),
  (x => 353, y => 164),
  (x => 354, y => 164),
  (x => 355, y => 164),
  (x => 366, y => 164),
  (x => 367, y => 164),
  (x => 368, y => 164),
  (x => 369, y => 164),
  (x => 370, y => 164),
  (x => 371, y => 164),
  (x => 372, y => 164),
  (x => 373, y => 164),
  (x => 249, y => 165),
  (x => 250, y => 165),
  (x => 251, y => 165),
  (x => 252, y => 165),
  (x => 253, y => 165),
  (x => 254, y => 165),
  (x => 255, y => 165),
  (x => 268, y => 165),
  (x => 269, y => 165),
  (x => 270, y => 165),
  (x => 271, y => 165),
  (x => 272, y => 165),
  (x => 273, y => 165),
  (x => 274, y => 165),
  (x => 275, y => 165),
  (x => 282, y => 165),
  (x => 283, y => 165),
  (x => 284, y => 165),
  (x => 285, y => 165),
  (x => 286, y => 165),
  (x => 287, y => 165),
  (x => 288, y => 165),
  (x => 289, y => 165),
  (x => 306, y => 165),
  (x => 307, y => 165),
  (x => 308, y => 165),
  (x => 309, y => 165),
  (x => 310, y => 165),
  (x => 311, y => 165),
  (x => 312, y => 165),
  (x => 313, y => 165),
  (x => 323, y => 165),
  (x => 324, y => 165),
  (x => 325, y => 165),
  (x => 326, y => 165),
  (x => 327, y => 165),
  (x => 328, y => 165),
  (x => 329, y => 165),
  (x => 332, y => 165),
  (x => 333, y => 165),
  (x => 334, y => 165),
  (x => 335, y => 165),
  (x => 336, y => 165),
  (x => 337, y => 165),
  (x => 349, y => 165),
  (x => 350, y => 165),
  (x => 351, y => 165),
  (x => 352, y => 165),
  (x => 353, y => 165),
  (x => 354, y => 165),
  (x => 355, y => 165),
  (x => 365, y => 165),
  (x => 366, y => 165),
  (x => 367, y => 165),
  (x => 368, y => 165),
  (x => 369, y => 165),
  (x => 370, y => 165),
  (x => 371, y => 165),
  (x => 372, y => 165),
  (x => 373, y => 165),
  (x => 249, y => 166),
  (x => 250, y => 166),
  (x => 251, y => 166),
  (x => 252, y => 166),
  (x => 253, y => 166),
  (x => 254, y => 166),
  (x => 255, y => 166),
  (x => 268, y => 166),
  (x => 269, y => 166),
  (x => 270, y => 166),
  (x => 271, y => 166),
  (x => 272, y => 166),
  (x => 273, y => 166),
  (x => 274, y => 166),
  (x => 275, y => 166),
  (x => 281, y => 166),
  (x => 282, y => 166),
  (x => 283, y => 166),
  (x => 284, y => 166),
  (x => 285, y => 166),
  (x => 286, y => 166),
  (x => 287, y => 166),
  (x => 288, y => 166),
  (x => 307, y => 166),
  (x => 308, y => 166),
  (x => 309, y => 166),
  (x => 310, y => 166),
  (x => 311, y => 166),
  (x => 312, y => 166),
  (x => 313, y => 166),
  (x => 314, y => 166),
  (x => 323, y => 166),
  (x => 324, y => 166),
  (x => 325, y => 166),
  (x => 326, y => 166),
  (x => 327, y => 166),
  (x => 328, y => 166),
  (x => 329, y => 166),
  (x => 332, y => 166),
  (x => 333, y => 166),
  (x => 334, y => 166),
  (x => 335, y => 166),
  (x => 336, y => 166),
  (x => 337, y => 166),
  (x => 338, y => 166),
  (x => 349, y => 166),
  (x => 350, y => 166),
  (x => 351, y => 166),
  (x => 352, y => 166),
  (x => 353, y => 166),
  (x => 354, y => 166),
  (x => 355, y => 166),
  (x => 365, y => 166),
  (x => 366, y => 166),
  (x => 367, y => 166),
  (x => 368, y => 166),
  (x => 369, y => 166),
  (x => 370, y => 166),
  (x => 371, y => 166),
  (x => 372, y => 166),
  (x => 249, y => 167),
  (x => 250, y => 167),
  (x => 251, y => 167),
  (x => 252, y => 167),
  (x => 253, y => 167),
  (x => 254, y => 167),
  (x => 255, y => 167),
  (x => 268, y => 167),
  (x => 269, y => 167),
  (x => 270, y => 167),
  (x => 271, y => 167),
  (x => 272, y => 167),
  (x => 273, y => 167),
  (x => 274, y => 167),
  (x => 275, y => 167),
  (x => 281, y => 167),
  (x => 282, y => 167),
  (x => 283, y => 167),
  (x => 284, y => 167),
  (x => 285, y => 167),
  (x => 286, y => 167),
  (x => 287, y => 167),
  (x => 288, y => 167),
  (x => 307, y => 167),
  (x => 308, y => 167),
  (x => 309, y => 167),
  (x => 310, y => 167),
  (x => 311, y => 167),
  (x => 312, y => 167),
  (x => 313, y => 167),
  (x => 314, y => 167),
  (x => 323, y => 167),
  (x => 324, y => 167),
  (x => 325, y => 167),
  (x => 326, y => 167),
  (x => 327, y => 167),
  (x => 328, y => 167),
  (x => 329, y => 167),
  (x => 332, y => 167),
  (x => 333, y => 167),
  (x => 334, y => 167),
  (x => 335, y => 167),
  (x => 336, y => 167),
  (x => 337, y => 167),
  (x => 338, y => 167),
  (x => 349, y => 167),
  (x => 350, y => 167),
  (x => 351, y => 167),
  (x => 352, y => 167),
  (x => 353, y => 167),
  (x => 354, y => 167),
  (x => 355, y => 167),
  (x => 365, y => 167),
  (x => 366, y => 167),
  (x => 367, y => 167),
  (x => 368, y => 167),
  (x => 369, y => 167),
  (x => 370, y => 167),
  (x => 371, y => 167),
  (x => 372, y => 167),
  (x => 249, y => 168),
  (x => 250, y => 168),
  (x => 251, y => 168),
  (x => 252, y => 168),
  (x => 253, y => 168),
  (x => 254, y => 168),
  (x => 255, y => 168),
  (x => 268, y => 168),
  (x => 269, y => 168),
  (x => 270, y => 168),
  (x => 271, y => 168),
  (x => 272, y => 168),
  (x => 273, y => 168),
  (x => 274, y => 168),
  (x => 275, y => 168),
  (x => 281, y => 168),
  (x => 282, y => 168),
  (x => 283, y => 168),
  (x => 284, y => 168),
  (x => 285, y => 168),
  (x => 286, y => 168),
  (x => 287, y => 168),
  (x => 307, y => 168),
  (x => 308, y => 168),
  (x => 309, y => 168),
  (x => 310, y => 168),
  (x => 311, y => 168),
  (x => 312, y => 168),
  (x => 313, y => 168),
  (x => 314, y => 168),
  (x => 323, y => 168),
  (x => 324, y => 168),
  (x => 325, y => 168),
  (x => 326, y => 168),
  (x => 327, y => 168),
  (x => 328, y => 168),
  (x => 329, y => 168),
  (x => 333, y => 168),
  (x => 334, y => 168),
  (x => 335, y => 168),
  (x => 336, y => 168),
  (x => 337, y => 168),
  (x => 338, y => 168),
  (x => 339, y => 168),
  (x => 349, y => 168),
  (x => 350, y => 168),
  (x => 351, y => 168),
  (x => 352, y => 168),
  (x => 353, y => 168),
  (x => 354, y => 168),
  (x => 355, y => 168),
  (x => 365, y => 168),
  (x => 366, y => 168),
  (x => 367, y => 168),
  (x => 368, y => 168),
  (x => 369, y => 168),
  (x => 370, y => 168),
  (x => 371, y => 168),
  (x => 249, y => 169),
  (x => 250, y => 169),
  (x => 251, y => 169),
  (x => 252, y => 169),
  (x => 253, y => 169),
  (x => 254, y => 169),
  (x => 255, y => 169),
  (x => 268, y => 169),
  (x => 269, y => 169),
  (x => 270, y => 169),
  (x => 271, y => 169),
  (x => 272, y => 169),
  (x => 273, y => 169),
  (x => 274, y => 169),
  (x => 281, y => 169),
  (x => 282, y => 169),
  (x => 283, y => 169),
  (x => 284, y => 169),
  (x => 285, y => 169),
  (x => 286, y => 169),
  (x => 287, y => 169),
  (x => 308, y => 169),
  (x => 309, y => 169),
  (x => 310, y => 169),
  (x => 311, y => 169),
  (x => 312, y => 169),
  (x => 313, y => 169),
  (x => 314, y => 169),
  (x => 323, y => 169),
  (x => 324, y => 169),
  (x => 325, y => 169),
  (x => 326, y => 169),
  (x => 327, y => 169),
  (x => 328, y => 169),
  (x => 329, y => 169),
  (x => 333, y => 169),
  (x => 334, y => 169),
  (x => 335, y => 169),
  (x => 336, y => 169),
  (x => 337, y => 169),
  (x => 338, y => 169),
  (x => 339, y => 169),
  (x => 349, y => 169),
  (x => 350, y => 169),
  (x => 351, y => 169),
  (x => 352, y => 169),
  (x => 353, y => 169),
  (x => 354, y => 169),
  (x => 355, y => 169),
  (x => 364, y => 169),
  (x => 365, y => 169),
  (x => 366, y => 169),
  (x => 367, y => 169),
  (x => 368, y => 169),
  (x => 369, y => 169),
  (x => 370, y => 169),
  (x => 371, y => 169),
  (x => 249, y => 170),
  (x => 250, y => 170),
  (x => 251, y => 170),
  (x => 252, y => 170),
  (x => 253, y => 170),
  (x => 254, y => 170),
  (x => 255, y => 170),
  (x => 268, y => 170),
  (x => 269, y => 170),
  (x => 270, y => 170),
  (x => 271, y => 170),
  (x => 272, y => 170),
  (x => 273, y => 170),
  (x => 274, y => 170),
  (x => 281, y => 170),
  (x => 282, y => 170),
  (x => 283, y => 170),
  (x => 284, y => 170),
  (x => 285, y => 170),
  (x => 286, y => 170),
  (x => 287, y => 170),
  (x => 308, y => 170),
  (x => 309, y => 170),
  (x => 310, y => 170),
  (x => 311, y => 170),
  (x => 312, y => 170),
  (x => 313, y => 170),
  (x => 314, y => 170),
  (x => 323, y => 170),
  (x => 324, y => 170),
  (x => 325, y => 170),
  (x => 326, y => 170),
  (x => 327, y => 170),
  (x => 328, y => 170),
  (x => 329, y => 170),
  (x => 334, y => 170),
  (x => 335, y => 170),
  (x => 336, y => 170),
  (x => 337, y => 170),
  (x => 338, y => 170),
  (x => 339, y => 170),
  (x => 340, y => 170),
  (x => 349, y => 170),
  (x => 350, y => 170),
  (x => 351, y => 170),
  (x => 352, y => 170),
  (x => 353, y => 170),
  (x => 354, y => 170),
  (x => 355, y => 170),
  (x => 364, y => 170),
  (x => 365, y => 170),
  (x => 366, y => 170),
  (x => 367, y => 170),
  (x => 368, y => 170),
  (x => 369, y => 170),
  (x => 370, y => 170),
  (x => 371, y => 170),
  (x => 249, y => 171),
  (x => 250, y => 171),
  (x => 251, y => 171),
  (x => 252, y => 171),
  (x => 253, y => 171),
  (x => 254, y => 171),
  (x => 255, y => 171),
  (x => 267, y => 171),
  (x => 268, y => 171),
  (x => 269, y => 171),
  (x => 270, y => 171),
  (x => 271, y => 171),
  (x => 272, y => 171),
  (x => 273, y => 171),
  (x => 274, y => 171),
  (x => 280, y => 171),
  (x => 281, y => 171),
  (x => 282, y => 171),
  (x => 283, y => 171),
  (x => 284, y => 171),
  (x => 285, y => 171),
  (x => 286, y => 171),
  (x => 287, y => 171),
  (x => 308, y => 171),
  (x => 309, y => 171),
  (x => 310, y => 171),
  (x => 311, y => 171),
  (x => 312, y => 171),
  (x => 313, y => 171),
  (x => 314, y => 171),
  (x => 323, y => 171),
  (x => 324, y => 171),
  (x => 325, y => 171),
  (x => 326, y => 171),
  (x => 327, y => 171),
  (x => 328, y => 171),
  (x => 329, y => 171),
  (x => 334, y => 171),
  (x => 335, y => 171),
  (x => 336, y => 171),
  (x => 337, y => 171),
  (x => 338, y => 171),
  (x => 339, y => 171),
  (x => 340, y => 171),
  (x => 349, y => 171),
  (x => 350, y => 171),
  (x => 351, y => 171),
  (x => 352, y => 171),
  (x => 353, y => 171),
  (x => 354, y => 171),
  (x => 355, y => 171),
  (x => 364, y => 171),
  (x => 365, y => 171),
  (x => 366, y => 171),
  (x => 367, y => 171),
  (x => 368, y => 171),
  (x => 369, y => 171),
  (x => 370, y => 171),
  (x => 371, y => 171),
  (x => 249, y => 172),
  (x => 250, y => 172),
  (x => 251, y => 172),
  (x => 252, y => 172),
  (x => 253, y => 172),
  (x => 254, y => 172),
  (x => 255, y => 172),
  (x => 267, y => 172),
  (x => 268, y => 172),
  (x => 269, y => 172),
  (x => 270, y => 172),
  (x => 271, y => 172),
  (x => 272, y => 172),
  (x => 273, y => 172),
  (x => 274, y => 172),
  (x => 280, y => 172),
  (x => 281, y => 172),
  (x => 282, y => 172),
  (x => 283, y => 172),
  (x => 284, y => 172),
  (x => 285, y => 172),
  (x => 286, y => 172),
  (x => 287, y => 172),
  (x => 308, y => 172),
  (x => 309, y => 172),
  (x => 310, y => 172),
  (x => 311, y => 172),
  (x => 312, y => 172),
  (x => 313, y => 172),
  (x => 314, y => 172),
  (x => 315, y => 172),
  (x => 323, y => 172),
  (x => 324, y => 172),
  (x => 325, y => 172),
  (x => 326, y => 172),
  (x => 327, y => 172),
  (x => 328, y => 172),
  (x => 329, y => 172),
  (x => 335, y => 172),
  (x => 336, y => 172),
  (x => 337, y => 172),
  (x => 338, y => 172),
  (x => 339, y => 172),
  (x => 340, y => 172),
  (x => 341, y => 172),
  (x => 349, y => 172),
  (x => 350, y => 172),
  (x => 351, y => 172),
  (x => 352, y => 172),
  (x => 353, y => 172),
  (x => 354, y => 172),
  (x => 355, y => 172),
  (x => 364, y => 172),
  (x => 365, y => 172),
  (x => 366, y => 172),
  (x => 367, y => 172),
  (x => 368, y => 172),
  (x => 369, y => 172),
  (x => 370, y => 172),
  (x => 371, y => 172),
  (x => 249, y => 173),
  (x => 250, y => 173),
  (x => 251, y => 173),
  (x => 252, y => 173),
  (x => 253, y => 173),
  (x => 254, y => 173),
  (x => 255, y => 173),
  (x => 266, y => 173),
  (x => 267, y => 173),
  (x => 268, y => 173),
  (x => 269, y => 173),
  (x => 270, y => 173),
  (x => 271, y => 173),
  (x => 272, y => 173),
  (x => 273, y => 173),
  (x => 274, y => 173),
  (x => 280, y => 173),
  (x => 281, y => 173),
  (x => 282, y => 173),
  (x => 283, y => 173),
  (x => 284, y => 173),
  (x => 285, y => 173),
  (x => 286, y => 173),
  (x => 287, y => 173),
  (x => 308, y => 173),
  (x => 309, y => 173),
  (x => 310, y => 173),
  (x => 311, y => 173),
  (x => 312, y => 173),
  (x => 313, y => 173),
  (x => 314, y => 173),
  (x => 315, y => 173),
  (x => 323, y => 173),
  (x => 324, y => 173),
  (x => 325, y => 173),
  (x => 326, y => 173),
  (x => 327, y => 173),
  (x => 328, y => 173),
  (x => 329, y => 173),
  (x => 335, y => 173),
  (x => 336, y => 173),
  (x => 337, y => 173),
  (x => 338, y => 173),
  (x => 339, y => 173),
  (x => 340, y => 173),
  (x => 341, y => 173),
  (x => 349, y => 173),
  (x => 350, y => 173),
  (x => 351, y => 173),
  (x => 352, y => 173),
  (x => 353, y => 173),
  (x => 354, y => 173),
  (x => 355, y => 173),
  (x => 364, y => 173),
  (x => 365, y => 173),
  (x => 366, y => 173),
  (x => 367, y => 173),
  (x => 368, y => 173),
  (x => 369, y => 173),
  (x => 370, y => 173),
  (x => 381, y => 173),
  (x => 382, y => 173),
  (x => 383, y => 173),
  (x => 384, y => 173),
  (x => 385, y => 173),
  (x => 386, y => 173),
  (x => 387, y => 173),
  (x => 388, y => 173),
  (x => 389, y => 173),
  (x => 390, y => 173),
  (x => 391, y => 173),
  (x => 392, y => 173),
  (x => 393, y => 173),
  (x => 394, y => 173),
  (x => 395, y => 173),
  (x => 249, y => 174),
  (x => 250, y => 174),
  (x => 251, y => 174),
  (x => 252, y => 174),
  (x => 253, y => 174),
  (x => 254, y => 174),
  (x => 255, y => 174),
  (x => 266, y => 174),
  (x => 267, y => 174),
  (x => 268, y => 174),
  (x => 269, y => 174),
  (x => 270, y => 174),
  (x => 271, y => 174),
  (x => 272, y => 174),
  (x => 273, y => 174),
  (x => 280, y => 174),
  (x => 281, y => 174),
  (x => 282, y => 174),
  (x => 283, y => 174),
  (x => 284, y => 174),
  (x => 285, y => 174),
  (x => 286, y => 174),
  (x => 287, y => 174),
  (x => 308, y => 174),
  (x => 309, y => 174),
  (x => 310, y => 174),
  (x => 311, y => 174),
  (x => 312, y => 174),
  (x => 313, y => 174),
  (x => 314, y => 174),
  (x => 315, y => 174),
  (x => 323, y => 174),
  (x => 324, y => 174),
  (x => 325, y => 174),
  (x => 326, y => 174),
  (x => 327, y => 174),
  (x => 328, y => 174),
  (x => 329, y => 174),
  (x => 336, y => 174),
  (x => 337, y => 174),
  (x => 338, y => 174),
  (x => 339, y => 174),
  (x => 340, y => 174),
  (x => 341, y => 174),
  (x => 342, y => 174),
  (x => 349, y => 174),
  (x => 350, y => 174),
  (x => 351, y => 174),
  (x => 352, y => 174),
  (x => 353, y => 174),
  (x => 354, y => 174),
  (x => 355, y => 174),
  (x => 364, y => 174),
  (x => 365, y => 174),
  (x => 366, y => 174),
  (x => 367, y => 174),
  (x => 368, y => 174),
  (x => 369, y => 174),
  (x => 370, y => 174),
  (x => 381, y => 174),
  (x => 382, y => 174),
  (x => 383, y => 174),
  (x => 384, y => 174),
  (x => 385, y => 174),
  (x => 386, y => 174),
  (x => 387, y => 174),
  (x => 388, y => 174),
  (x => 389, y => 174),
  (x => 390, y => 174),
  (x => 391, y => 174),
  (x => 392, y => 174),
  (x => 393, y => 174),
  (x => 394, y => 174),
  (x => 395, y => 174),
  (x => 249, y => 175),
  (x => 250, y => 175),
  (x => 251, y => 175),
  (x => 252, y => 175),
  (x => 253, y => 175),
  (x => 254, y => 175),
  (x => 255, y => 175),
  (x => 256, y => 175),
  (x => 264, y => 175),
  (x => 265, y => 175),
  (x => 266, y => 175),
  (x => 267, y => 175),
  (x => 268, y => 175),
  (x => 269, y => 175),
  (x => 270, y => 175),
  (x => 271, y => 175),
  (x => 272, y => 175),
  (x => 273, y => 175),
  (x => 280, y => 175),
  (x => 281, y => 175),
  (x => 282, y => 175),
  (x => 283, y => 175),
  (x => 284, y => 175),
  (x => 285, y => 175),
  (x => 286, y => 175),
  (x => 287, y => 175),
  (x => 308, y => 175),
  (x => 309, y => 175),
  (x => 310, y => 175),
  (x => 311, y => 175),
  (x => 312, y => 175),
  (x => 313, y => 175),
  (x => 314, y => 175),
  (x => 315, y => 175),
  (x => 323, y => 175),
  (x => 324, y => 175),
  (x => 325, y => 175),
  (x => 326, y => 175),
  (x => 327, y => 175),
  (x => 328, y => 175),
  (x => 329, y => 175),
  (x => 336, y => 175),
  (x => 337, y => 175),
  (x => 338, y => 175),
  (x => 339, y => 175),
  (x => 340, y => 175),
  (x => 341, y => 175),
  (x => 342, y => 175),
  (x => 349, y => 175),
  (x => 350, y => 175),
  (x => 351, y => 175),
  (x => 352, y => 175),
  (x => 353, y => 175),
  (x => 354, y => 175),
  (x => 355, y => 175),
  (x => 364, y => 175),
  (x => 365, y => 175),
  (x => 366, y => 175),
  (x => 367, y => 175),
  (x => 368, y => 175),
  (x => 369, y => 175),
  (x => 370, y => 175),
  (x => 381, y => 175),
  (x => 382, y => 175),
  (x => 383, y => 175),
  (x => 384, y => 175),
  (x => 385, y => 175),
  (x => 386, y => 175),
  (x => 387, y => 175),
  (x => 388, y => 175),
  (x => 389, y => 175),
  (x => 390, y => 175),
  (x => 391, y => 175),
  (x => 392, y => 175),
  (x => 393, y => 175),
  (x => 394, y => 175),
  (x => 395, y => 175),
  (x => 249, y => 176),
  (x => 250, y => 176),
  (x => 251, y => 176),
  (x => 252, y => 176),
  (x => 253, y => 176),
  (x => 254, y => 176),
  (x => 255, y => 176),
  (x => 256, y => 176),
  (x => 257, y => 176),
  (x => 258, y => 176),
  (x => 259, y => 176),
  (x => 260, y => 176),
  (x => 261, y => 176),
  (x => 262, y => 176),
  (x => 263, y => 176),
  (x => 264, y => 176),
  (x => 265, y => 176),
  (x => 266, y => 176),
  (x => 267, y => 176),
  (x => 268, y => 176),
  (x => 269, y => 176),
  (x => 270, y => 176),
  (x => 271, y => 176),
  (x => 272, y => 176),
  (x => 280, y => 176),
  (x => 281, y => 176),
  (x => 282, y => 176),
  (x => 283, y => 176),
  (x => 284, y => 176),
  (x => 285, y => 176),
  (x => 286, y => 176),
  (x => 287, y => 176),
  (x => 308, y => 176),
  (x => 309, y => 176),
  (x => 310, y => 176),
  (x => 311, y => 176),
  (x => 312, y => 176),
  (x => 313, y => 176),
  (x => 314, y => 176),
  (x => 315, y => 176),
  (x => 323, y => 176),
  (x => 324, y => 176),
  (x => 325, y => 176),
  (x => 326, y => 176),
  (x => 327, y => 176),
  (x => 328, y => 176),
  (x => 329, y => 176),
  (x => 337, y => 176),
  (x => 338, y => 176),
  (x => 339, y => 176),
  (x => 340, y => 176),
  (x => 341, y => 176),
  (x => 342, y => 176),
  (x => 343, y => 176),
  (x => 349, y => 176),
  (x => 350, y => 176),
  (x => 351, y => 176),
  (x => 352, y => 176),
  (x => 353, y => 176),
  (x => 354, y => 176),
  (x => 355, y => 176),
  (x => 364, y => 176),
  (x => 365, y => 176),
  (x => 366, y => 176),
  (x => 367, y => 176),
  (x => 368, y => 176),
  (x => 369, y => 176),
  (x => 370, y => 176),
  (x => 381, y => 176),
  (x => 382, y => 176),
  (x => 383, y => 176),
  (x => 384, y => 176),
  (x => 385, y => 176),
  (x => 386, y => 176),
  (x => 387, y => 176),
  (x => 388, y => 176),
  (x => 389, y => 176),
  (x => 390, y => 176),
  (x => 391, y => 176),
  (x => 392, y => 176),
  (x => 393, y => 176),
  (x => 394, y => 176),
  (x => 395, y => 176),
  (x => 249, y => 177),
  (x => 250, y => 177),
  (x => 251, y => 177),
  (x => 252, y => 177),
  (x => 253, y => 177),
  (x => 254, y => 177),
  (x => 255, y => 177),
  (x => 256, y => 177),
  (x => 257, y => 177),
  (x => 258, y => 177),
  (x => 259, y => 177),
  (x => 260, y => 177),
  (x => 261, y => 177),
  (x => 262, y => 177),
  (x => 263, y => 177),
  (x => 264, y => 177),
  (x => 265, y => 177),
  (x => 266, y => 177),
  (x => 267, y => 177),
  (x => 268, y => 177),
  (x => 269, y => 177),
  (x => 270, y => 177),
  (x => 271, y => 177),
  (x => 272, y => 177),
  (x => 280, y => 177),
  (x => 281, y => 177),
  (x => 282, y => 177),
  (x => 283, y => 177),
  (x => 284, y => 177),
  (x => 285, y => 177),
  (x => 286, y => 177),
  (x => 287, y => 177),
  (x => 308, y => 177),
  (x => 309, y => 177),
  (x => 310, y => 177),
  (x => 311, y => 177),
  (x => 312, y => 177),
  (x => 313, y => 177),
  (x => 314, y => 177),
  (x => 315, y => 177),
  (x => 323, y => 177),
  (x => 324, y => 177),
  (x => 325, y => 177),
  (x => 326, y => 177),
  (x => 327, y => 177),
  (x => 328, y => 177),
  (x => 329, y => 177),
  (x => 337, y => 177),
  (x => 338, y => 177),
  (x => 339, y => 177),
  (x => 340, y => 177),
  (x => 341, y => 177),
  (x => 342, y => 177),
  (x => 343, y => 177),
  (x => 349, y => 177),
  (x => 350, y => 177),
  (x => 351, y => 177),
  (x => 352, y => 177),
  (x => 353, y => 177),
  (x => 354, y => 177),
  (x => 355, y => 177),
  (x => 364, y => 177),
  (x => 365, y => 177),
  (x => 366, y => 177),
  (x => 367, y => 177),
  (x => 368, y => 177),
  (x => 369, y => 177),
  (x => 370, y => 177),
  (x => 381, y => 177),
  (x => 382, y => 177),
  (x => 383, y => 177),
  (x => 384, y => 177),
  (x => 385, y => 177),
  (x => 386, y => 177),
  (x => 387, y => 177),
  (x => 388, y => 177),
  (x => 389, y => 177),
  (x => 390, y => 177),
  (x => 391, y => 177),
  (x => 392, y => 177),
  (x => 393, y => 177),
  (x => 394, y => 177),
  (x => 395, y => 177),
  (x => 249, y => 178),
  (x => 250, y => 178),
  (x => 251, y => 178),
  (x => 252, y => 178),
  (x => 253, y => 178),
  (x => 254, y => 178),
  (x => 255, y => 178),
  (x => 256, y => 178),
  (x => 257, y => 178),
  (x => 258, y => 178),
  (x => 259, y => 178),
  (x => 260, y => 178),
  (x => 261, y => 178),
  (x => 262, y => 178),
  (x => 263, y => 178),
  (x => 264, y => 178),
  (x => 265, y => 178),
  (x => 266, y => 178),
  (x => 267, y => 178),
  (x => 268, y => 178),
  (x => 269, y => 178),
  (x => 270, y => 178),
  (x => 271, y => 178),
  (x => 280, y => 178),
  (x => 281, y => 178),
  (x => 282, y => 178),
  (x => 283, y => 178),
  (x => 284, y => 178),
  (x => 285, y => 178),
  (x => 286, y => 178),
  (x => 287, y => 178),
  (x => 308, y => 178),
  (x => 309, y => 178),
  (x => 310, y => 178),
  (x => 311, y => 178),
  (x => 312, y => 178),
  (x => 313, y => 178),
  (x => 314, y => 178),
  (x => 315, y => 178),
  (x => 323, y => 178),
  (x => 324, y => 178),
  (x => 325, y => 178),
  (x => 326, y => 178),
  (x => 327, y => 178),
  (x => 328, y => 178),
  (x => 329, y => 178),
  (x => 338, y => 178),
  (x => 339, y => 178),
  (x => 340, y => 178),
  (x => 341, y => 178),
  (x => 342, y => 178),
  (x => 343, y => 178),
  (x => 344, y => 178),
  (x => 349, y => 178),
  (x => 350, y => 178),
  (x => 351, y => 178),
  (x => 352, y => 178),
  (x => 353, y => 178),
  (x => 354, y => 178),
  (x => 355, y => 178),
  (x => 364, y => 178),
  (x => 365, y => 178),
  (x => 366, y => 178),
  (x => 367, y => 178),
  (x => 368, y => 178),
  (x => 369, y => 178),
  (x => 370, y => 178),
  (x => 381, y => 178),
  (x => 382, y => 178),
  (x => 383, y => 178),
  (x => 384, y => 178),
  (x => 385, y => 178),
  (x => 386, y => 178),
  (x => 387, y => 178),
  (x => 388, y => 178),
  (x => 389, y => 178),
  (x => 390, y => 178),
  (x => 391, y => 178),
  (x => 392, y => 178),
  (x => 393, y => 178),
  (x => 394, y => 178),
  (x => 395, y => 178),
  (x => 249, y => 179),
  (x => 250, y => 179),
  (x => 251, y => 179),
  (x => 252, y => 179),
  (x => 253, y => 179),
  (x => 254, y => 179),
  (x => 255, y => 179),
  (x => 256, y => 179),
  (x => 257, y => 179),
  (x => 258, y => 179),
  (x => 259, y => 179),
  (x => 260, y => 179),
  (x => 261, y => 179),
  (x => 262, y => 179),
  (x => 263, y => 179),
  (x => 264, y => 179),
  (x => 265, y => 179),
  (x => 266, y => 179),
  (x => 267, y => 179),
  (x => 268, y => 179),
  (x => 269, y => 179),
  (x => 270, y => 179),
  (x => 280, y => 179),
  (x => 281, y => 179),
  (x => 282, y => 179),
  (x => 283, y => 179),
  (x => 284, y => 179),
  (x => 285, y => 179),
  (x => 286, y => 179),
  (x => 287, y => 179),
  (x => 308, y => 179),
  (x => 309, y => 179),
  (x => 310, y => 179),
  (x => 311, y => 179),
  (x => 312, y => 179),
  (x => 313, y => 179),
  (x => 314, y => 179),
  (x => 315, y => 179),
  (x => 323, y => 179),
  (x => 324, y => 179),
  (x => 325, y => 179),
  (x => 326, y => 179),
  (x => 327, y => 179),
  (x => 328, y => 179),
  (x => 329, y => 179),
  (x => 338, y => 179),
  (x => 339, y => 179),
  (x => 340, y => 179),
  (x => 341, y => 179),
  (x => 342, y => 179),
  (x => 343, y => 179),
  (x => 344, y => 179),
  (x => 349, y => 179),
  (x => 350, y => 179),
  (x => 351, y => 179),
  (x => 352, y => 179),
  (x => 353, y => 179),
  (x => 354, y => 179),
  (x => 355, y => 179),
  (x => 364, y => 179),
  (x => 365, y => 179),
  (x => 366, y => 179),
  (x => 367, y => 179),
  (x => 368, y => 179),
  (x => 369, y => 179),
  (x => 370, y => 179),
  (x => 381, y => 179),
  (x => 382, y => 179),
  (x => 383, y => 179),
  (x => 384, y => 179),
  (x => 385, y => 179),
  (x => 386, y => 179),
  (x => 387, y => 179),
  (x => 388, y => 179),
  (x => 389, y => 179),
  (x => 390, y => 179),
  (x => 391, y => 179),
  (x => 392, y => 179),
  (x => 393, y => 179),
  (x => 394, y => 179),
  (x => 395, y => 179),
  (x => 249, y => 180),
  (x => 250, y => 180),
  (x => 251, y => 180),
  (x => 252, y => 180),
  (x => 253, y => 180),
  (x => 254, y => 180),
  (x => 255, y => 180),
  (x => 256, y => 180),
  (x => 257, y => 180),
  (x => 258, y => 180),
  (x => 259, y => 180),
  (x => 260, y => 180),
  (x => 261, y => 180),
  (x => 262, y => 180),
  (x => 263, y => 180),
  (x => 264, y => 180),
  (x => 265, y => 180),
  (x => 266, y => 180),
  (x => 267, y => 180),
  (x => 268, y => 180),
  (x => 269, y => 180),
  (x => 280, y => 180),
  (x => 281, y => 180),
  (x => 282, y => 180),
  (x => 283, y => 180),
  (x => 284, y => 180),
  (x => 285, y => 180),
  (x => 286, y => 180),
  (x => 287, y => 180),
  (x => 308, y => 180),
  (x => 309, y => 180),
  (x => 310, y => 180),
  (x => 311, y => 180),
  (x => 312, y => 180),
  (x => 313, y => 180),
  (x => 314, y => 180),
  (x => 323, y => 180),
  (x => 324, y => 180),
  (x => 325, y => 180),
  (x => 326, y => 180),
  (x => 327, y => 180),
  (x => 328, y => 180),
  (x => 329, y => 180),
  (x => 339, y => 180),
  (x => 340, y => 180),
  (x => 341, y => 180),
  (x => 342, y => 180),
  (x => 343, y => 180),
  (x => 344, y => 180),
  (x => 349, y => 180),
  (x => 350, y => 180),
  (x => 351, y => 180),
  (x => 352, y => 180),
  (x => 353, y => 180),
  (x => 354, y => 180),
  (x => 355, y => 180),
  (x => 364, y => 180),
  (x => 365, y => 180),
  (x => 366, y => 180),
  (x => 367, y => 180),
  (x => 368, y => 180),
  (x => 369, y => 180),
  (x => 370, y => 180),
  (x => 381, y => 180),
  (x => 382, y => 180),
  (x => 383, y => 180),
  (x => 384, y => 180),
  (x => 385, y => 180),
  (x => 386, y => 180),
  (x => 387, y => 180),
  (x => 388, y => 180),
  (x => 389, y => 180),
  (x => 390, y => 180),
  (x => 391, y => 180),
  (x => 392, y => 180),
  (x => 393, y => 180),
  (x => 394, y => 180),
  (x => 395, y => 180),
  (x => 249, y => 181),
  (x => 250, y => 181),
  (x => 251, y => 181),
  (x => 252, y => 181),
  (x => 253, y => 181),
  (x => 254, y => 181),
  (x => 255, y => 181),
  (x => 256, y => 181),
  (x => 257, y => 181),
  (x => 258, y => 181),
  (x => 259, y => 181),
  (x => 260, y => 181),
  (x => 261, y => 181),
  (x => 262, y => 181),
  (x => 263, y => 181),
  (x => 264, y => 181),
  (x => 265, y => 181),
  (x => 266, y => 181),
  (x => 267, y => 181),
  (x => 268, y => 181),
  (x => 280, y => 181),
  (x => 281, y => 181),
  (x => 282, y => 181),
  (x => 283, y => 181),
  (x => 284, y => 181),
  (x => 285, y => 181),
  (x => 286, y => 181),
  (x => 287, y => 181),
  (x => 308, y => 181),
  (x => 309, y => 181),
  (x => 310, y => 181),
  (x => 311, y => 181),
  (x => 312, y => 181),
  (x => 313, y => 181),
  (x => 314, y => 181),
  (x => 323, y => 181),
  (x => 324, y => 181),
  (x => 325, y => 181),
  (x => 326, y => 181),
  (x => 327, y => 181),
  (x => 328, y => 181),
  (x => 329, y => 181),
  (x => 339, y => 181),
  (x => 340, y => 181),
  (x => 341, y => 181),
  (x => 342, y => 181),
  (x => 343, y => 181),
  (x => 344, y => 181),
  (x => 345, y => 181),
  (x => 349, y => 181),
  (x => 350, y => 181),
  (x => 351, y => 181),
  (x => 352, y => 181),
  (x => 353, y => 181),
  (x => 354, y => 181),
  (x => 355, y => 181),
  (x => 364, y => 181),
  (x => 365, y => 181),
  (x => 366, y => 181),
  (x => 367, y => 181),
  (x => 368, y => 181),
  (x => 369, y => 181),
  (x => 370, y => 181),
  (x => 371, y => 181),
  (x => 389, y => 181),
  (x => 390, y => 181),
  (x => 391, y => 181),
  (x => 392, y => 181),
  (x => 393, y => 181),
  (x => 394, y => 181),
  (x => 395, y => 181),
  (x => 249, y => 182),
  (x => 250, y => 182),
  (x => 251, y => 182),
  (x => 252, y => 182),
  (x => 253, y => 182),
  (x => 254, y => 182),
  (x => 255, y => 182),
  (x => 256, y => 182),
  (x => 257, y => 182),
  (x => 258, y => 182),
  (x => 259, y => 182),
  (x => 260, y => 182),
  (x => 261, y => 182),
  (x => 262, y => 182),
  (x => 263, y => 182),
  (x => 264, y => 182),
  (x => 265, y => 182),
  (x => 280, y => 182),
  (x => 281, y => 182),
  (x => 282, y => 182),
  (x => 283, y => 182),
  (x => 284, y => 182),
  (x => 285, y => 182),
  (x => 286, y => 182),
  (x => 287, y => 182),
  (x => 308, y => 182),
  (x => 309, y => 182),
  (x => 310, y => 182),
  (x => 311, y => 182),
  (x => 312, y => 182),
  (x => 313, y => 182),
  (x => 314, y => 182),
  (x => 323, y => 182),
  (x => 324, y => 182),
  (x => 325, y => 182),
  (x => 326, y => 182),
  (x => 327, y => 182),
  (x => 328, y => 182),
  (x => 329, y => 182),
  (x => 340, y => 182),
  (x => 341, y => 182),
  (x => 342, y => 182),
  (x => 343, y => 182),
  (x => 344, y => 182),
  (x => 345, y => 182),
  (x => 346, y => 182),
  (x => 350, y => 182),
  (x => 351, y => 182),
  (x => 352, y => 182),
  (x => 353, y => 182),
  (x => 354, y => 182),
  (x => 355, y => 182),
  (x => 364, y => 182),
  (x => 365, y => 182),
  (x => 366, y => 182),
  (x => 367, y => 182),
  (x => 368, y => 182),
  (x => 369, y => 182),
  (x => 370, y => 182),
  (x => 371, y => 182),
  (x => 389, y => 182),
  (x => 390, y => 182),
  (x => 391, y => 182),
  (x => 392, y => 182),
  (x => 393, y => 182),
  (x => 394, y => 182),
  (x => 395, y => 182),
  (x => 249, y => 183),
  (x => 250, y => 183),
  (x => 251, y => 183),
  (x => 252, y => 183),
  (x => 253, y => 183),
  (x => 254, y => 183),
  (x => 255, y => 183),
  (x => 256, y => 183),
  (x => 281, y => 183),
  (x => 282, y => 183),
  (x => 283, y => 183),
  (x => 284, y => 183),
  (x => 285, y => 183),
  (x => 286, y => 183),
  (x => 287, y => 183),
  (x => 307, y => 183),
  (x => 308, y => 183),
  (x => 309, y => 183),
  (x => 310, y => 183),
  (x => 311, y => 183),
  (x => 312, y => 183),
  (x => 313, y => 183),
  (x => 314, y => 183),
  (x => 323, y => 183),
  (x => 324, y => 183),
  (x => 325, y => 183),
  (x => 326, y => 183),
  (x => 327, y => 183),
  (x => 328, y => 183),
  (x => 329, y => 183),
  (x => 340, y => 183),
  (x => 341, y => 183),
  (x => 342, y => 183),
  (x => 343, y => 183),
  (x => 344, y => 183),
  (x => 345, y => 183),
  (x => 346, y => 183),
  (x => 350, y => 183),
  (x => 351, y => 183),
  (x => 352, y => 183),
  (x => 353, y => 183),
  (x => 354, y => 183),
  (x => 355, y => 183),
  (x => 364, y => 183),
  (x => 365, y => 183),
  (x => 366, y => 183),
  (x => 367, y => 183),
  (x => 368, y => 183),
  (x => 369, y => 183),
  (x => 370, y => 183),
  (x => 371, y => 183),
  (x => 389, y => 183),
  (x => 390, y => 183),
  (x => 391, y => 183),
  (x => 392, y => 183),
  (x => 393, y => 183),
  (x => 394, y => 183),
  (x => 395, y => 183),
  (x => 249, y => 184),
  (x => 250, y => 184),
  (x => 251, y => 184),
  (x => 252, y => 184),
  (x => 253, y => 184),
  (x => 254, y => 184),
  (x => 255, y => 184),
  (x => 281, y => 184),
  (x => 282, y => 184),
  (x => 283, y => 184),
  (x => 284, y => 184),
  (x => 285, y => 184),
  (x => 286, y => 184),
  (x => 287, y => 184),
  (x => 288, y => 184),
  (x => 307, y => 184),
  (x => 308, y => 184),
  (x => 309, y => 184),
  (x => 310, y => 184),
  (x => 311, y => 184),
  (x => 312, y => 184),
  (x => 313, y => 184),
  (x => 314, y => 184),
  (x => 323, y => 184),
  (x => 324, y => 184),
  (x => 325, y => 184),
  (x => 326, y => 184),
  (x => 327, y => 184),
  (x => 328, y => 184),
  (x => 329, y => 184),
  (x => 341, y => 184),
  (x => 342, y => 184),
  (x => 343, y => 184),
  (x => 344, y => 184),
  (x => 345, y => 184),
  (x => 346, y => 184),
  (x => 350, y => 184),
  (x => 351, y => 184),
  (x => 352, y => 184),
  (x => 353, y => 184),
  (x => 354, y => 184),
  (x => 355, y => 184),
  (x => 364, y => 184),
  (x => 365, y => 184),
  (x => 366, y => 184),
  (x => 367, y => 184),
  (x => 368, y => 184),
  (x => 369, y => 184),
  (x => 370, y => 184),
  (x => 371, y => 184),
  (x => 389, y => 184),
  (x => 390, y => 184),
  (x => 391, y => 184),
  (x => 392, y => 184),
  (x => 393, y => 184),
  (x => 394, y => 184),
  (x => 395, y => 184),
  (x => 249, y => 185),
  (x => 250, y => 185),
  (x => 251, y => 185),
  (x => 252, y => 185),
  (x => 253, y => 185),
  (x => 254, y => 185),
  (x => 255, y => 185),
  (x => 281, y => 185),
  (x => 282, y => 185),
  (x => 283, y => 185),
  (x => 284, y => 185),
  (x => 285, y => 185),
  (x => 286, y => 185),
  (x => 287, y => 185),
  (x => 288, y => 185),
  (x => 307, y => 185),
  (x => 308, y => 185),
  (x => 309, y => 185),
  (x => 310, y => 185),
  (x => 311, y => 185),
  (x => 312, y => 185),
  (x => 313, y => 185),
  (x => 314, y => 185),
  (x => 323, y => 185),
  (x => 324, y => 185),
  (x => 325, y => 185),
  (x => 326, y => 185),
  (x => 327, y => 185),
  (x => 328, y => 185),
  (x => 329, y => 185),
  (x => 341, y => 185),
  (x => 342, y => 185),
  (x => 343, y => 185),
  (x => 344, y => 185),
  (x => 345, y => 185),
  (x => 346, y => 185),
  (x => 347, y => 185),
  (x => 350, y => 185),
  (x => 351, y => 185),
  (x => 352, y => 185),
  (x => 353, y => 185),
  (x => 354, y => 185),
  (x => 355, y => 185),
  (x => 365, y => 185),
  (x => 366, y => 185),
  (x => 367, y => 185),
  (x => 368, y => 185),
  (x => 369, y => 185),
  (x => 370, y => 185),
  (x => 371, y => 185),
  (x => 372, y => 185),
  (x => 389, y => 185),
  (x => 390, y => 185),
  (x => 391, y => 185),
  (x => 392, y => 185),
  (x => 393, y => 185),
  (x => 394, y => 185),
  (x => 395, y => 185),
  (x => 249, y => 186),
  (x => 250, y => 186),
  (x => 251, y => 186),
  (x => 252, y => 186),
  (x => 253, y => 186),
  (x => 254, y => 186),
  (x => 255, y => 186),
  (x => 281, y => 186),
  (x => 282, y => 186),
  (x => 283, y => 186),
  (x => 284, y => 186),
  (x => 285, y => 186),
  (x => 286, y => 186),
  (x => 287, y => 186),
  (x => 288, y => 186),
  (x => 307, y => 186),
  (x => 308, y => 186),
  (x => 309, y => 186),
  (x => 310, y => 186),
  (x => 311, y => 186),
  (x => 312, y => 186),
  (x => 313, y => 186),
  (x => 323, y => 186),
  (x => 324, y => 186),
  (x => 325, y => 186),
  (x => 326, y => 186),
  (x => 327, y => 186),
  (x => 328, y => 186),
  (x => 329, y => 186),
  (x => 342, y => 186),
  (x => 343, y => 186),
  (x => 344, y => 186),
  (x => 345, y => 186),
  (x => 346, y => 186),
  (x => 347, y => 186),
  (x => 348, y => 186),
  (x => 349, y => 186),
  (x => 350, y => 186),
  (x => 351, y => 186),
  (x => 352, y => 186),
  (x => 353, y => 186),
  (x => 354, y => 186),
  (x => 355, y => 186),
  (x => 365, y => 186),
  (x => 366, y => 186),
  (x => 367, y => 186),
  (x => 368, y => 186),
  (x => 369, y => 186),
  (x => 370, y => 186),
  (x => 371, y => 186),
  (x => 372, y => 186),
  (x => 389, y => 186),
  (x => 390, y => 186),
  (x => 391, y => 186),
  (x => 392, y => 186),
  (x => 393, y => 186),
  (x => 394, y => 186),
  (x => 395, y => 186),
  (x => 249, y => 187),
  (x => 250, y => 187),
  (x => 251, y => 187),
  (x => 252, y => 187),
  (x => 253, y => 187),
  (x => 254, y => 187),
  (x => 255, y => 187),
  (x => 281, y => 187),
  (x => 282, y => 187),
  (x => 283, y => 187),
  (x => 284, y => 187),
  (x => 285, y => 187),
  (x => 286, y => 187),
  (x => 287, y => 187),
  (x => 288, y => 187),
  (x => 289, y => 187),
  (x => 306, y => 187),
  (x => 307, y => 187),
  (x => 308, y => 187),
  (x => 309, y => 187),
  (x => 310, y => 187),
  (x => 311, y => 187),
  (x => 312, y => 187),
  (x => 313, y => 187),
  (x => 323, y => 187),
  (x => 324, y => 187),
  (x => 325, y => 187),
  (x => 326, y => 187),
  (x => 327, y => 187),
  (x => 328, y => 187),
  (x => 329, y => 187),
  (x => 342, y => 187),
  (x => 343, y => 187),
  (x => 344, y => 187),
  (x => 345, y => 187),
  (x => 346, y => 187),
  (x => 347, y => 187),
  (x => 348, y => 187),
  (x => 349, y => 187),
  (x => 350, y => 187),
  (x => 351, y => 187),
  (x => 352, y => 187),
  (x => 353, y => 187),
  (x => 354, y => 187),
  (x => 355, y => 187),
  (x => 365, y => 187),
  (x => 366, y => 187),
  (x => 367, y => 187),
  (x => 368, y => 187),
  (x => 369, y => 187),
  (x => 370, y => 187),
  (x => 371, y => 187),
  (x => 372, y => 187),
  (x => 389, y => 187),
  (x => 390, y => 187),
  (x => 391, y => 187),
  (x => 392, y => 187),
  (x => 393, y => 187),
  (x => 394, y => 187),
  (x => 395, y => 187),
  (x => 249, y => 188),
  (x => 250, y => 188),
  (x => 251, y => 188),
  (x => 252, y => 188),
  (x => 253, y => 188),
  (x => 254, y => 188),
  (x => 255, y => 188),
  (x => 282, y => 188),
  (x => 283, y => 188),
  (x => 284, y => 188),
  (x => 285, y => 188),
  (x => 286, y => 188),
  (x => 287, y => 188),
  (x => 288, y => 188),
  (x => 289, y => 188),
  (x => 306, y => 188),
  (x => 307, y => 188),
  (x => 308, y => 188),
  (x => 309, y => 188),
  (x => 310, y => 188),
  (x => 311, y => 188),
  (x => 312, y => 188),
  (x => 313, y => 188),
  (x => 323, y => 188),
  (x => 324, y => 188),
  (x => 325, y => 188),
  (x => 326, y => 188),
  (x => 327, y => 188),
  (x => 328, y => 188),
  (x => 329, y => 188),
  (x => 343, y => 188),
  (x => 344, y => 188),
  (x => 345, y => 188),
  (x => 346, y => 188),
  (x => 347, y => 188),
  (x => 348, y => 188),
  (x => 349, y => 188),
  (x => 350, y => 188),
  (x => 351, y => 188),
  (x => 352, y => 188),
  (x => 353, y => 188),
  (x => 354, y => 188),
  (x => 355, y => 188),
  (x => 365, y => 188),
  (x => 366, y => 188),
  (x => 367, y => 188),
  (x => 368, y => 188),
  (x => 369, y => 188),
  (x => 370, y => 188),
  (x => 371, y => 188),
  (x => 372, y => 188),
  (x => 373, y => 188),
  (x => 389, y => 188),
  (x => 390, y => 188),
  (x => 391, y => 188),
  (x => 392, y => 188),
  (x => 393, y => 188),
  (x => 394, y => 188),
  (x => 395, y => 188),
  (x => 249, y => 189),
  (x => 250, y => 189),
  (x => 251, y => 189),
  (x => 252, y => 189),
  (x => 253, y => 189),
  (x => 254, y => 189),
  (x => 255, y => 189),
  (x => 282, y => 189),
  (x => 283, y => 189),
  (x => 284, y => 189),
  (x => 285, y => 189),
  (x => 286, y => 189),
  (x => 287, y => 189),
  (x => 288, y => 189),
  (x => 289, y => 189),
  (x => 290, y => 189),
  (x => 305, y => 189),
  (x => 306, y => 189),
  (x => 307, y => 189),
  (x => 308, y => 189),
  (x => 309, y => 189),
  (x => 310, y => 189),
  (x => 311, y => 189),
  (x => 312, y => 189),
  (x => 323, y => 189),
  (x => 324, y => 189),
  (x => 325, y => 189),
  (x => 326, y => 189),
  (x => 327, y => 189),
  (x => 328, y => 189),
  (x => 329, y => 189),
  (x => 343, y => 189),
  (x => 344, y => 189),
  (x => 345, y => 189),
  (x => 346, y => 189),
  (x => 347, y => 189),
  (x => 348, y => 189),
  (x => 349, y => 189),
  (x => 350, y => 189),
  (x => 351, y => 189),
  (x => 352, y => 189),
  (x => 353, y => 189),
  (x => 354, y => 189),
  (x => 355, y => 189),
  (x => 366, y => 189),
  (x => 367, y => 189),
  (x => 368, y => 189),
  (x => 369, y => 189),
  (x => 370, y => 189),
  (x => 371, y => 189),
  (x => 372, y => 189),
  (x => 373, y => 189),
  (x => 374, y => 189),
  (x => 389, y => 189),
  (x => 390, y => 189),
  (x => 391, y => 189),
  (x => 392, y => 189),
  (x => 393, y => 189),
  (x => 394, y => 189),
  (x => 395, y => 189),
  (x => 249, y => 190),
  (x => 250, y => 190),
  (x => 251, y => 190),
  (x => 252, y => 190),
  (x => 253, y => 190),
  (x => 254, y => 190),
  (x => 255, y => 190),
  (x => 283, y => 190),
  (x => 284, y => 190),
  (x => 285, y => 190),
  (x => 286, y => 190),
  (x => 287, y => 190),
  (x => 288, y => 190),
  (x => 289, y => 190),
  (x => 290, y => 190),
  (x => 291, y => 190),
  (x => 304, y => 190),
  (x => 305, y => 190),
  (x => 306, y => 190),
  (x => 307, y => 190),
  (x => 308, y => 190),
  (x => 309, y => 190),
  (x => 310, y => 190),
  (x => 311, y => 190),
  (x => 312, y => 190),
  (x => 323, y => 190),
  (x => 324, y => 190),
  (x => 325, y => 190),
  (x => 326, y => 190),
  (x => 327, y => 190),
  (x => 328, y => 190),
  (x => 329, y => 190),
  (x => 344, y => 190),
  (x => 345, y => 190),
  (x => 346, y => 190),
  (x => 347, y => 190),
  (x => 348, y => 190),
  (x => 349, y => 190),
  (x => 350, y => 190),
  (x => 351, y => 190),
  (x => 352, y => 190),
  (x => 353, y => 190),
  (x => 354, y => 190),
  (x => 355, y => 190),
  (x => 366, y => 190),
  (x => 367, y => 190),
  (x => 368, y => 190),
  (x => 369, y => 190),
  (x => 370, y => 190),
  (x => 371, y => 190),
  (x => 372, y => 190),
  (x => 373, y => 190),
  (x => 374, y => 190),
  (x => 375, y => 190),
  (x => 389, y => 190),
  (x => 390, y => 190),
  (x => 391, y => 190),
  (x => 392, y => 190),
  (x => 393, y => 190),
  (x => 394, y => 190),
  (x => 395, y => 190),
  (x => 249, y => 191),
  (x => 250, y => 191),
  (x => 251, y => 191),
  (x => 252, y => 191),
  (x => 253, y => 191),
  (x => 254, y => 191),
  (x => 255, y => 191),
  (x => 283, y => 191),
  (x => 284, y => 191),
  (x => 285, y => 191),
  (x => 286, y => 191),
  (x => 287, y => 191),
  (x => 288, y => 191),
  (x => 289, y => 191),
  (x => 290, y => 191),
  (x => 291, y => 191),
  (x => 292, y => 191),
  (x => 303, y => 191),
  (x => 304, y => 191),
  (x => 305, y => 191),
  (x => 306, y => 191),
  (x => 307, y => 191),
  (x => 308, y => 191),
  (x => 309, y => 191),
  (x => 310, y => 191),
  (x => 311, y => 191),
  (x => 312, y => 191),
  (x => 323, y => 191),
  (x => 324, y => 191),
  (x => 325, y => 191),
  (x => 326, y => 191),
  (x => 327, y => 191),
  (x => 328, y => 191),
  (x => 329, y => 191),
  (x => 344, y => 191),
  (x => 345, y => 191),
  (x => 346, y => 191),
  (x => 347, y => 191),
  (x => 348, y => 191),
  (x => 349, y => 191),
  (x => 350, y => 191),
  (x => 351, y => 191),
  (x => 352, y => 191),
  (x => 353, y => 191),
  (x => 354, y => 191),
  (x => 355, y => 191),
  (x => 367, y => 191),
  (x => 368, y => 191),
  (x => 369, y => 191),
  (x => 370, y => 191),
  (x => 371, y => 191),
  (x => 372, y => 191),
  (x => 373, y => 191),
  (x => 374, y => 191),
  (x => 375, y => 191),
  (x => 376, y => 191),
  (x => 389, y => 191),
  (x => 390, y => 191),
  (x => 391, y => 191),
  (x => 392, y => 191),
  (x => 393, y => 191),
  (x => 394, y => 191),
  (x => 395, y => 191),
  (x => 249, y => 192),
  (x => 250, y => 192),
  (x => 251, y => 192),
  (x => 252, y => 192),
  (x => 253, y => 192),
  (x => 254, y => 192),
  (x => 255, y => 192),
  (x => 284, y => 192),
  (x => 285, y => 192),
  (x => 286, y => 192),
  (x => 287, y => 192),
  (x => 288, y => 192),
  (x => 289, y => 192),
  (x => 290, y => 192),
  (x => 291, y => 192),
  (x => 292, y => 192),
  (x => 293, y => 192),
  (x => 301, y => 192),
  (x => 302, y => 192),
  (x => 303, y => 192),
  (x => 304, y => 192),
  (x => 305, y => 192),
  (x => 306, y => 192),
  (x => 307, y => 192),
  (x => 308, y => 192),
  (x => 309, y => 192),
  (x => 310, y => 192),
  (x => 311, y => 192),
  (x => 323, y => 192),
  (x => 324, y => 192),
  (x => 325, y => 192),
  (x => 326, y => 192),
  (x => 327, y => 192),
  (x => 328, y => 192),
  (x => 329, y => 192),
  (x => 345, y => 192),
  (x => 346, y => 192),
  (x => 347, y => 192),
  (x => 348, y => 192),
  (x => 349, y => 192),
  (x => 350, y => 192),
  (x => 351, y => 192),
  (x => 352, y => 192),
  (x => 353, y => 192),
  (x => 354, y => 192),
  (x => 355, y => 192),
  (x => 367, y => 192),
  (x => 368, y => 192),
  (x => 369, y => 192),
  (x => 370, y => 192),
  (x => 371, y => 192),
  (x => 372, y => 192),
  (x => 373, y => 192),
  (x => 374, y => 192),
  (x => 375, y => 192),
  (x => 376, y => 192),
  (x => 377, y => 192),
  (x => 388, y => 192),
  (x => 389, y => 192),
  (x => 390, y => 192),
  (x => 391, y => 192),
  (x => 392, y => 192),
  (x => 393, y => 192),
  (x => 394, y => 192),
  (x => 395, y => 192),
  (x => 249, y => 193),
  (x => 250, y => 193),
  (x => 251, y => 193),
  (x => 252, y => 193),
  (x => 253, y => 193),
  (x => 254, y => 193),
  (x => 255, y => 193),
  (x => 284, y => 193),
  (x => 285, y => 193),
  (x => 286, y => 193),
  (x => 287, y => 193),
  (x => 288, y => 193),
  (x => 289, y => 193),
  (x => 290, y => 193),
  (x => 291, y => 193),
  (x => 292, y => 193),
  (x => 293, y => 193),
  (x => 294, y => 193),
  (x => 295, y => 193),
  (x => 296, y => 193),
  (x => 297, y => 193),
  (x => 298, y => 193),
  (x => 299, y => 193),
  (x => 300, y => 193),
  (x => 301, y => 193),
  (x => 302, y => 193),
  (x => 303, y => 193),
  (x => 304, y => 193),
  (x => 305, y => 193),
  (x => 306, y => 193),
  (x => 307, y => 193),
  (x => 308, y => 193),
  (x => 309, y => 193),
  (x => 310, y => 193),
  (x => 323, y => 193),
  (x => 324, y => 193),
  (x => 325, y => 193),
  (x => 326, y => 193),
  (x => 327, y => 193),
  (x => 328, y => 193),
  (x => 329, y => 193),
  (x => 345, y => 193),
  (x => 346, y => 193),
  (x => 347, y => 193),
  (x => 348, y => 193),
  (x => 349, y => 193),
  (x => 350, y => 193),
  (x => 351, y => 193),
  (x => 352, y => 193),
  (x => 353, y => 193),
  (x => 354, y => 193),
  (x => 355, y => 193),
  (x => 368, y => 193),
  (x => 369, y => 193),
  (x => 370, y => 193),
  (x => 371, y => 193),
  (x => 372, y => 193),
  (x => 373, y => 193),
  (x => 374, y => 193),
  (x => 375, y => 193),
  (x => 376, y => 193),
  (x => 377, y => 193),
  (x => 378, y => 193),
  (x => 379, y => 193),
  (x => 380, y => 193),
  (x => 381, y => 193),
  (x => 385, y => 193),
  (x => 386, y => 193),
  (x => 387, y => 193),
  (x => 388, y => 193),
  (x => 389, y => 193),
  (x => 390, y => 193),
  (x => 391, y => 193),
  (x => 392, y => 193),
  (x => 393, y => 193),
  (x => 394, y => 193),
  (x => 395, y => 193),
  (x => 249, y => 194),
  (x => 250, y => 194),
  (x => 251, y => 194),
  (x => 252, y => 194),
  (x => 253, y => 194),
  (x => 254, y => 194),
  (x => 255, y => 194),
  (x => 285, y => 194),
  (x => 286, y => 194),
  (x => 287, y => 194),
  (x => 288, y => 194),
  (x => 289, y => 194),
  (x => 290, y => 194),
  (x => 291, y => 194),
  (x => 292, y => 194),
  (x => 293, y => 194),
  (x => 294, y => 194),
  (x => 295, y => 194),
  (x => 296, y => 194),
  (x => 297, y => 194),
  (x => 298, y => 194),
  (x => 299, y => 194),
  (x => 300, y => 194),
  (x => 301, y => 194),
  (x => 302, y => 194),
  (x => 303, y => 194),
  (x => 304, y => 194),
  (x => 305, y => 194),
  (x => 306, y => 194),
  (x => 307, y => 194),
  (x => 308, y => 194),
  (x => 309, y => 194),
  (x => 310, y => 194),
  (x => 323, y => 194),
  (x => 324, y => 194),
  (x => 325, y => 194),
  (x => 326, y => 194),
  (x => 327, y => 194),
  (x => 328, y => 194),
  (x => 329, y => 194),
  (x => 346, y => 194),
  (x => 347, y => 194),
  (x => 348, y => 194),
  (x => 349, y => 194),
  (x => 350, y => 194),
  (x => 351, y => 194),
  (x => 352, y => 194),
  (x => 353, y => 194),
  (x => 354, y => 194),
  (x => 355, y => 194),
  (x => 368, y => 194),
  (x => 369, y => 194),
  (x => 370, y => 194),
  (x => 371, y => 194),
  (x => 372, y => 194),
  (x => 373, y => 194),
  (x => 374, y => 194),
  (x => 375, y => 194),
  (x => 376, y => 194),
  (x => 377, y => 194),
  (x => 378, y => 194),
  (x => 379, y => 194),
  (x => 380, y => 194),
  (x => 381, y => 194),
  (x => 382, y => 194),
  (x => 383, y => 194),
  (x => 384, y => 194),
  (x => 385, y => 194),
  (x => 386, y => 194),
  (x => 387, y => 194),
  (x => 388, y => 194),
  (x => 389, y => 194),
  (x => 390, y => 194),
  (x => 391, y => 194),
  (x => 392, y => 194),
  (x => 393, y => 194),
  (x => 394, y => 194),
  (x => 395, y => 194),
  (x => 249, y => 195),
  (x => 250, y => 195),
  (x => 251, y => 195),
  (x => 252, y => 195),
  (x => 253, y => 195),
  (x => 254, y => 195),
  (x => 255, y => 195),
  (x => 285, y => 195),
  (x => 286, y => 195),
  (x => 287, y => 195),
  (x => 288, y => 195),
  (x => 289, y => 195),
  (x => 290, y => 195),
  (x => 291, y => 195),
  (x => 292, y => 195),
  (x => 293, y => 195),
  (x => 294, y => 195),
  (x => 295, y => 195),
  (x => 296, y => 195),
  (x => 297, y => 195),
  (x => 298, y => 195),
  (x => 299, y => 195),
  (x => 300, y => 195),
  (x => 301, y => 195),
  (x => 302, y => 195),
  (x => 303, y => 195),
  (x => 304, y => 195),
  (x => 305, y => 195),
  (x => 306, y => 195),
  (x => 307, y => 195),
  (x => 308, y => 195),
  (x => 309, y => 195),
  (x => 323, y => 195),
  (x => 324, y => 195),
  (x => 325, y => 195),
  (x => 326, y => 195),
  (x => 327, y => 195),
  (x => 328, y => 195),
  (x => 329, y => 195),
  (x => 346, y => 195),
  (x => 347, y => 195),
  (x => 348, y => 195),
  (x => 349, y => 195),
  (x => 350, y => 195),
  (x => 351, y => 195),
  (x => 352, y => 195),
  (x => 353, y => 195),
  (x => 354, y => 195),
  (x => 355, y => 195),
  (x => 369, y => 195),
  (x => 370, y => 195),
  (x => 371, y => 195),
  (x => 372, y => 195),
  (x => 373, y => 195),
  (x => 374, y => 195),
  (x => 375, y => 195),
  (x => 376, y => 195),
  (x => 377, y => 195),
  (x => 378, y => 195),
  (x => 379, y => 195),
  (x => 380, y => 195),
  (x => 381, y => 195),
  (x => 382, y => 195),
  (x => 383, y => 195),
  (x => 384, y => 195),
  (x => 385, y => 195),
  (x => 386, y => 195),
  (x => 387, y => 195),
  (x => 388, y => 195),
  (x => 389, y => 195),
  (x => 390, y => 195),
  (x => 391, y => 195),
  (x => 392, y => 195),
  (x => 393, y => 195),
  (x => 394, y => 195),
  (x => 395, y => 195),
  (x => 249, y => 196),
  (x => 250, y => 196),
  (x => 251, y => 196),
  (x => 252, y => 196),
  (x => 253, y => 196),
  (x => 254, y => 196),
  (x => 255, y => 196),
  (x => 286, y => 196),
  (x => 287, y => 196),
  (x => 288, y => 196),
  (x => 289, y => 196),
  (x => 290, y => 196),
  (x => 291, y => 196),
  (x => 292, y => 196),
  (x => 293, y => 196),
  (x => 294, y => 196),
  (x => 295, y => 196),
  (x => 296, y => 196),
  (x => 297, y => 196),
  (x => 298, y => 196),
  (x => 299, y => 196),
  (x => 300, y => 196),
  (x => 301, y => 196),
  (x => 302, y => 196),
  (x => 303, y => 196),
  (x => 304, y => 196),
  (x => 305, y => 196),
  (x => 306, y => 196),
  (x => 307, y => 196),
  (x => 308, y => 196),
  (x => 323, y => 196),
  (x => 324, y => 196),
  (x => 325, y => 196),
  (x => 326, y => 196),
  (x => 327, y => 196),
  (x => 328, y => 196),
  (x => 329, y => 196),
  (x => 347, y => 196),
  (x => 348, y => 196),
  (x => 349, y => 196),
  (x => 350, y => 196),
  (x => 351, y => 196),
  (x => 352, y => 196),
  (x => 353, y => 196),
  (x => 354, y => 196),
  (x => 355, y => 196),
  (x => 370, y => 196),
  (x => 371, y => 196),
  (x => 372, y => 196),
  (x => 373, y => 196),
  (x => 374, y => 196),
  (x => 375, y => 196),
  (x => 376, y => 196),
  (x => 377, y => 196),
  (x => 378, y => 196),
  (x => 379, y => 196),
  (x => 380, y => 196),
  (x => 381, y => 196),
  (x => 382, y => 196),
  (x => 383, y => 196),
  (x => 384, y => 196),
  (x => 385, y => 196),
  (x => 386, y => 196),
  (x => 387, y => 196),
  (x => 388, y => 196),
  (x => 389, y => 196),
  (x => 390, y => 196),
  (x => 391, y => 196),
  (x => 392, y => 196),
  (x => 393, y => 196),
  (x => 394, y => 196),
  (x => 395, y => 196),
  (x => 249, y => 197),
  (x => 250, y => 197),
  (x => 251, y => 197),
  (x => 252, y => 197),
  (x => 253, y => 197),
  (x => 254, y => 197),
  (x => 255, y => 197),
  (x => 287, y => 197),
  (x => 288, y => 197),
  (x => 289, y => 197),
  (x => 290, y => 197),
  (x => 291, y => 197),
  (x => 292, y => 197),
  (x => 293, y => 197),
  (x => 294, y => 197),
  (x => 295, y => 197),
  (x => 296, y => 197),
  (x => 297, y => 197),
  (x => 298, y => 197),
  (x => 299, y => 197),
  (x => 300, y => 197),
  (x => 301, y => 197),
  (x => 302, y => 197),
  (x => 303, y => 197),
  (x => 304, y => 197),
  (x => 305, y => 197),
  (x => 306, y => 197),
  (x => 307, y => 197),
  (x => 323, y => 197),
  (x => 324, y => 197),
  (x => 325, y => 197),
  (x => 326, y => 197),
  (x => 327, y => 197),
  (x => 328, y => 197),
  (x => 329, y => 197),
  (x => 347, y => 197),
  (x => 348, y => 197),
  (x => 349, y => 197),
  (x => 350, y => 197),
  (x => 351, y => 197),
  (x => 352, y => 197),
  (x => 353, y => 197),
  (x => 354, y => 197),
  (x => 355, y => 197),
  (x => 371, y => 197),
  (x => 372, y => 197),
  (x => 373, y => 197),
  (x => 374, y => 197),
  (x => 375, y => 197),
  (x => 376, y => 197),
  (x => 377, y => 197),
  (x => 378, y => 197),
  (x => 379, y => 197),
  (x => 380, y => 197),
  (x => 381, y => 197),
  (x => 382, y => 197),
  (x => 383, y => 197),
  (x => 384, y => 197),
  (x => 385, y => 197),
  (x => 386, y => 197),
  (x => 387, y => 197),
  (x => 388, y => 197),
  (x => 389, y => 197),
  (x => 390, y => 197),
  (x => 391, y => 197),
  (x => 392, y => 197),
  (x => 393, y => 197),
  (x => 394, y => 197),
  (x => 395, y => 197),
  (x => 249, y => 198),
  (x => 250, y => 198),
  (x => 251, y => 198),
  (x => 252, y => 198),
  (x => 253, y => 198),
  (x => 254, y => 198),
  (x => 255, y => 198),
  (x => 288, y => 198),
  (x => 289, y => 198),
  (x => 290, y => 198),
  (x => 291, y => 198),
  (x => 292, y => 198),
  (x => 293, y => 198),
  (x => 294, y => 198),
  (x => 295, y => 198),
  (x => 296, y => 198),
  (x => 297, y => 198),
  (x => 298, y => 198),
  (x => 299, y => 198),
  (x => 300, y => 198),
  (x => 301, y => 198),
  (x => 302, y => 198),
  (x => 303, y => 198),
  (x => 304, y => 198),
  (x => 305, y => 198),
  (x => 306, y => 198),
  (x => 323, y => 198),
  (x => 324, y => 198),
  (x => 325, y => 198),
  (x => 326, y => 198),
  (x => 327, y => 198),
  (x => 328, y => 198),
  (x => 329, y => 198),
  (x => 348, y => 198),
  (x => 349, y => 198),
  (x => 350, y => 198),
  (x => 351, y => 198),
  (x => 352, y => 198),
  (x => 353, y => 198),
  (x => 354, y => 198),
  (x => 355, y => 198),
  (x => 372, y => 198),
  (x => 373, y => 198),
  (x => 374, y => 198),
  (x => 375, y => 198),
  (x => 376, y => 198),
  (x => 377, y => 198),
  (x => 378, y => 198),
  (x => 379, y => 198),
  (x => 380, y => 198),
  (x => 381, y => 198),
  (x => 382, y => 198),
  (x => 383, y => 198),
  (x => 384, y => 198),
  (x => 385, y => 198),
  (x => 386, y => 198),
  (x => 387, y => 198),
  (x => 388, y => 198),
  (x => 389, y => 198),
  (x => 390, y => 198),
  (x => 391, y => 198),
  (x => 392, y => 198),
  (x => 393, y => 198),
  (x => 394, y => 198),
  (x => 249, y => 199),
  (x => 250, y => 199),
  (x => 251, y => 199),
  (x => 252, y => 199),
  (x => 253, y => 199),
  (x => 254, y => 199),
  (x => 255, y => 199),
  (x => 290, y => 199),
  (x => 291, y => 199),
  (x => 292, y => 199),
  (x => 293, y => 199),
  (x => 294, y => 199),
  (x => 295, y => 199),
  (x => 296, y => 199),
  (x => 297, y => 199),
  (x => 298, y => 199),
  (x => 299, y => 199),
  (x => 300, y => 199),
  (x => 301, y => 199),
  (x => 302, y => 199),
  (x => 303, y => 199),
  (x => 304, y => 199),
  (x => 305, y => 199),
  (x => 323, y => 199),
  (x => 324, y => 199),
  (x => 325, y => 199),
  (x => 326, y => 199),
  (x => 327, y => 199),
  (x => 328, y => 199),
  (x => 329, y => 199),
  (x => 348, y => 199),
  (x => 349, y => 199),
  (x => 350, y => 199),
  (x => 351, y => 199),
  (x => 352, y => 199),
  (x => 353, y => 199),
  (x => 354, y => 199),
  (x => 355, y => 199),
  (x => 374, y => 199),
  (x => 375, y => 199),
  (x => 376, y => 199),
  (x => 377, y => 199),
  (x => 378, y => 199),
  (x => 379, y => 199),
  (x => 380, y => 199),
  (x => 381, y => 199),
  (x => 382, y => 199),
  (x => 383, y => 199),
  (x => 384, y => 199),
  (x => 385, y => 199),
  (x => 386, y => 199),
  (x => 387, y => 199),
  (x => 388, y => 199),
  (x => 389, y => 199),
  (x => 390, y => 199),
  (x => 391, y => 199),
  (x => 392, y => 199),
  (x => 249, y => 200),
  (x => 250, y => 200),
  (x => 251, y => 200),
  (x => 252, y => 200),
  (x => 253, y => 200),
  (x => 254, y => 200),
  (x => 255, y => 200),
  (x => 256, y => 200),
  (x => 292, y => 200),
  (x => 293, y => 200),
  (x => 294, y => 200),
  (x => 295, y => 200),
  (x => 296, y => 200),
  (x => 297, y => 200),
  (x => 298, y => 200),
  (x => 299, y => 200),
  (x => 300, y => 200),
  (x => 301, y => 200),
  (x => 302, y => 200),
  (x => 303, y => 200),
  (x => 323, y => 200),
  (x => 324, y => 200),
  (x => 325, y => 200),
  (x => 326, y => 200),
  (x => 327, y => 200),
  (x => 328, y => 200),
  (x => 329, y => 200),
  (x => 348, y => 200),
  (x => 349, y => 200),
  (x => 350, y => 200),
  (x => 351, y => 200),
  (x => 352, y => 200),
  (x => 353, y => 200),
  (x => 354, y => 200),
  (x => 355, y => 200),
  (x => 376, y => 200),
  (x => 377, y => 200),
  (x => 378, y => 200),
  (x => 379, y => 200),
  (x => 380, y => 200),
  (x => 381, y => 200),
  (x => 382, y => 200),
  (x => 383, y => 200),
  (x => 384, y => 200),
  (x => 385, y => 200),
  (x => 386, y => 200),
  (x => 387, y => 200),
  (x => 388, y => 200),
  (x => 389, y => 200),
  (x => 295, y => 201),
  (x => 296, y => 201),
  (x => 297, y => 201),
  (x => 298, y => 201),
  (x => 299, y => 201),
  (x => 380, y => 201),
  (x => 381, y => 201),
  (x => 382, y => 201),
  (x => 383, y => 201),
  (x => 384, y => 201),
  (x => 385, y => 201),
  (x => 377, y => 255),
  (x => 378, y => 255),
  (x => 265, y => 256),
  (x => 266, y => 256),
  (x => 267, y => 256),
  (x => 268, y => 256),
  (x => 269, y => 256),
  (x => 270, y => 256),
  (x => 271, y => 256),
  (x => 272, y => 256),
  (x => 273, y => 256),
  (x => 274, y => 256),
  (x => 275, y => 256),
  (x => 350, y => 256),
  (x => 351, y => 256),
  (x => 352, y => 256),
  (x => 353, y => 256),
  (x => 354, y => 256),
  (x => 355, y => 256),
  (x => 356, y => 256),
  (x => 357, y => 256),
  (x => 358, y => 256),
  (x => 359, y => 256),
  (x => 360, y => 256),
  (x => 376, y => 256),
  (x => 377, y => 256),
  (x => 378, y => 256),
  (x => 265, y => 257),
  (x => 266, y => 257),
  (x => 267, y => 257),
  (x => 268, y => 257),
  (x => 269, y => 257),
  (x => 270, y => 257),
  (x => 271, y => 257),
  (x => 272, y => 257),
  (x => 273, y => 257),
  (x => 274, y => 257),
  (x => 275, y => 257),
  (x => 276, y => 257),
  (x => 350, y => 257),
  (x => 351, y => 257),
  (x => 352, y => 257),
  (x => 353, y => 257),
  (x => 354, y => 257),
  (x => 355, y => 257),
  (x => 356, y => 257),
  (x => 357, y => 257),
  (x => 358, y => 257),
  (x => 359, y => 257),
  (x => 360, y => 257),
  (x => 361, y => 257),
  (x => 362, y => 257),
  (x => 375, y => 257),
  (x => 376, y => 257),
  (x => 377, y => 257),
  (x => 378, y => 257),
  (x => 265, y => 258),
  (x => 266, y => 258),
  (x => 267, y => 258),
  (x => 268, y => 258),
  (x => 269, y => 258),
  (x => 270, y => 258),
  (x => 271, y => 258),
  (x => 272, y => 258),
  (x => 273, y => 258),
  (x => 274, y => 258),
  (x => 275, y => 258),
  (x => 276, y => 258),
  (x => 277, y => 258),
  (x => 350, y => 258),
  (x => 351, y => 258),
  (x => 352, y => 258),
  (x => 353, y => 258),
  (x => 354, y => 258),
  (x => 355, y => 258),
  (x => 356, y => 258),
  (x => 357, y => 258),
  (x => 358, y => 258),
  (x => 359, y => 258),
  (x => 360, y => 258),
  (x => 361, y => 258),
  (x => 362, y => 258),
  (x => 373, y => 258),
  (x => 374, y => 258),
  (x => 375, y => 258),
  (x => 376, y => 258),
  (x => 377, y => 258),
  (x => 378, y => 258),
  (x => 265, y => 259),
  (x => 266, y => 259),
  (x => 267, y => 259),
  (x => 268, y => 259),
  (x => 269, y => 259),
  (x => 270, y => 259),
  (x => 271, y => 259),
  (x => 272, y => 259),
  (x => 273, y => 259),
  (x => 274, y => 259),
  (x => 275, y => 259),
  (x => 276, y => 259),
  (x => 277, y => 259),
  (x => 278, y => 259),
  (x => 350, y => 259),
  (x => 351, y => 259),
  (x => 352, y => 259),
  (x => 353, y => 259),
  (x => 357, y => 259),
  (x => 358, y => 259),
  (x => 359, y => 259),
  (x => 360, y => 259),
  (x => 361, y => 259),
  (x => 362, y => 259),
  (x => 363, y => 259),
  (x => 371, y => 259),
  (x => 372, y => 259),
  (x => 373, y => 259),
  (x => 374, y => 259),
  (x => 375, y => 259),
  (x => 376, y => 259),
  (x => 377, y => 259),
  (x => 378, y => 259),
  (x => 265, y => 260),
  (x => 266, y => 260),
  (x => 267, y => 260),
  (x => 268, y => 260),
  (x => 274, y => 260),
  (x => 275, y => 260),
  (x => 276, y => 260),
  (x => 277, y => 260),
  (x => 278, y => 260),
  (x => 350, y => 260),
  (x => 351, y => 260),
  (x => 352, y => 260),
  (x => 353, y => 260),
  (x => 360, y => 260),
  (x => 361, y => 260),
  (x => 362, y => 260),
  (x => 363, y => 260),
  (x => 371, y => 260),
  (x => 372, y => 260),
  (x => 373, y => 260),
  (x => 374, y => 260),
  (x => 375, y => 260),
  (x => 376, y => 260),
  (x => 377, y => 260),
  (x => 378, y => 260),
  (x => 265, y => 261),
  (x => 266, y => 261),
  (x => 267, y => 261),
  (x => 268, y => 261),
  (x => 275, y => 261),
  (x => 276, y => 261),
  (x => 277, y => 261),
  (x => 278, y => 261),
  (x => 350, y => 261),
  (x => 351, y => 261),
  (x => 352, y => 261),
  (x => 353, y => 261),
  (x => 360, y => 261),
  (x => 361, y => 261),
  (x => 362, y => 261),
  (x => 363, y => 261),
  (x => 371, y => 261),
  (x => 372, y => 261),
  (x => 373, y => 261),
  (x => 374, y => 261),
  (x => 375, y => 261),
  (x => 376, y => 261),
  (x => 377, y => 261),
  (x => 378, y => 261),
  (x => 265, y => 262),
  (x => 266, y => 262),
  (x => 267, y => 262),
  (x => 268, y => 262),
  (x => 276, y => 262),
  (x => 277, y => 262),
  (x => 278, y => 262),
  (x => 279, y => 262),
  (x => 350, y => 262),
  (x => 351, y => 262),
  (x => 352, y => 262),
  (x => 353, y => 262),
  (x => 361, y => 262),
  (x => 362, y => 262),
  (x => 363, y => 262),
  (x => 371, y => 262),
  (x => 372, y => 262),
  (x => 373, y => 262),
  (x => 376, y => 262),
  (x => 377, y => 262),
  (x => 378, y => 262),
  (x => 265, y => 263),
  (x => 266, y => 263),
  (x => 267, y => 263),
  (x => 268, y => 263),
  (x => 276, y => 263),
  (x => 277, y => 263),
  (x => 278, y => 263),
  (x => 279, y => 263),
  (x => 350, y => 263),
  (x => 351, y => 263),
  (x => 352, y => 263),
  (x => 353, y => 263),
  (x => 361, y => 263),
  (x => 362, y => 263),
  (x => 363, y => 263),
  (x => 371, y => 263),
  (x => 376, y => 263),
  (x => 377, y => 263),
  (x => 378, y => 263),
  (x => 265, y => 264),
  (x => 266, y => 264),
  (x => 267, y => 264),
  (x => 268, y => 264),
  (x => 276, y => 264),
  (x => 277, y => 264),
  (x => 278, y => 264),
  (x => 279, y => 264),
  (x => 284, y => 264),
  (x => 285, y => 264),
  (x => 286, y => 264),
  (x => 290, y => 264),
  (x => 291, y => 264),
  (x => 292, y => 264),
  (x => 300, y => 264),
  (x => 301, y => 264),
  (x => 302, y => 264),
  (x => 303, y => 264),
  (x => 304, y => 264),
  (x => 315, y => 264),
  (x => 316, y => 264),
  (x => 317, y => 264),
  (x => 318, y => 264),
  (x => 319, y => 264),
  (x => 320, y => 264),
  (x => 321, y => 264),
  (x => 329, y => 264),
  (x => 330, y => 264),
  (x => 331, y => 264),
  (x => 332, y => 264),
  (x => 333, y => 264),
  (x => 334, y => 264),
  (x => 335, y => 264),
  (x => 350, y => 264),
  (x => 351, y => 264),
  (x => 352, y => 264),
  (x => 353, y => 264),
  (x => 361, y => 264),
  (x => 362, y => 264),
  (x => 363, y => 264),
  (x => 376, y => 264),
  (x => 377, y => 264),
  (x => 378, y => 264),
  (x => 265, y => 265),
  (x => 266, y => 265),
  (x => 267, y => 265),
  (x => 268, y => 265),
  (x => 276, y => 265),
  (x => 277, y => 265),
  (x => 278, y => 265),
  (x => 279, y => 265),
  (x => 284, y => 265),
  (x => 285, y => 265),
  (x => 286, y => 265),
  (x => 290, y => 265),
  (x => 291, y => 265),
  (x => 292, y => 265),
  (x => 298, y => 265),
  (x => 299, y => 265),
  (x => 300, y => 265),
  (x => 301, y => 265),
  (x => 302, y => 265),
  (x => 303, y => 265),
  (x => 304, y => 265),
  (x => 305, y => 265),
  (x => 306, y => 265),
  (x => 314, y => 265),
  (x => 315, y => 265),
  (x => 316, y => 265),
  (x => 317, y => 265),
  (x => 318, y => 265),
  (x => 319, y => 265),
  (x => 320, y => 265),
  (x => 321, y => 265),
  (x => 328, y => 265),
  (x => 329, y => 265),
  (x => 330, y => 265),
  (x => 331, y => 265),
  (x => 332, y => 265),
  (x => 333, y => 265),
  (x => 334, y => 265),
  (x => 335, y => 265),
  (x => 350, y => 265),
  (x => 351, y => 265),
  (x => 352, y => 265),
  (x => 353, y => 265),
  (x => 360, y => 265),
  (x => 361, y => 265),
  (x => 362, y => 265),
  (x => 363, y => 265),
  (x => 376, y => 265),
  (x => 377, y => 265),
  (x => 378, y => 265),
  (x => 265, y => 266),
  (x => 266, y => 266),
  (x => 267, y => 266),
  (x => 268, y => 266),
  (x => 276, y => 266),
  (x => 277, y => 266),
  (x => 278, y => 266),
  (x => 279, y => 266),
  (x => 284, y => 266),
  (x => 285, y => 266),
  (x => 286, y => 266),
  (x => 289, y => 266),
  (x => 290, y => 266),
  (x => 291, y => 266),
  (x => 292, y => 266),
  (x => 298, y => 266),
  (x => 299, y => 266),
  (x => 300, y => 266),
  (x => 301, y => 266),
  (x => 302, y => 266),
  (x => 303, y => 266),
  (x => 304, y => 266),
  (x => 305, y => 266),
  (x => 306, y => 266),
  (x => 313, y => 266),
  (x => 314, y => 266),
  (x => 315, y => 266),
  (x => 316, y => 266),
  (x => 317, y => 266),
  (x => 318, y => 266),
  (x => 319, y => 266),
  (x => 320, y => 266),
  (x => 321, y => 266),
  (x => 327, y => 266),
  (x => 328, y => 266),
  (x => 329, y => 266),
  (x => 330, y => 266),
  (x => 331, y => 266),
  (x => 332, y => 266),
  (x => 333, y => 266),
  (x => 334, y => 266),
  (x => 335, y => 266),
  (x => 350, y => 266),
  (x => 351, y => 266),
  (x => 352, y => 266),
  (x => 353, y => 266),
  (x => 360, y => 266),
  (x => 361, y => 266),
  (x => 362, y => 266),
  (x => 376, y => 266),
  (x => 377, y => 266),
  (x => 378, y => 266),
  (x => 265, y => 267),
  (x => 266, y => 267),
  (x => 267, y => 267),
  (x => 268, y => 267),
  (x => 276, y => 267),
  (x => 277, y => 267),
  (x => 278, y => 267),
  (x => 284, y => 267),
  (x => 285, y => 267),
  (x => 286, y => 267),
  (x => 289, y => 267),
  (x => 290, y => 267),
  (x => 291, y => 267),
  (x => 292, y => 267),
  (x => 297, y => 267),
  (x => 298, y => 267),
  (x => 299, y => 267),
  (x => 300, y => 267),
  (x => 304, y => 267),
  (x => 305, y => 267),
  (x => 306, y => 267),
  (x => 307, y => 267),
  (x => 313, y => 267),
  (x => 314, y => 267),
  (x => 315, y => 267),
  (x => 321, y => 267),
  (x => 326, y => 267),
  (x => 327, y => 267),
  (x => 328, y => 267),
  (x => 329, y => 267),
  (x => 335, y => 267),
  (x => 350, y => 267),
  (x => 351, y => 267),
  (x => 352, y => 267),
  (x => 353, y => 267),
  (x => 358, y => 267),
  (x => 359, y => 267),
  (x => 360, y => 267),
  (x => 361, y => 267),
  (x => 376, y => 267),
  (x => 377, y => 267),
  (x => 378, y => 267),
  (x => 265, y => 268),
  (x => 266, y => 268),
  (x => 267, y => 268),
  (x => 268, y => 268),
  (x => 275, y => 268),
  (x => 276, y => 268),
  (x => 277, y => 268),
  (x => 278, y => 268),
  (x => 284, y => 268),
  (x => 285, y => 268),
  (x => 286, y => 268),
  (x => 287, y => 268),
  (x => 288, y => 268),
  (x => 289, y => 268),
  (x => 296, y => 268),
  (x => 297, y => 268),
  (x => 298, y => 268),
  (x => 299, y => 268),
  (x => 305, y => 268),
  (x => 306, y => 268),
  (x => 307, y => 268),
  (x => 312, y => 268),
  (x => 313, y => 268),
  (x => 314, y => 268),
  (x => 315, y => 268),
  (x => 326, y => 268),
  (x => 327, y => 268),
  (x => 328, y => 268),
  (x => 350, y => 268),
  (x => 351, y => 268),
  (x => 352, y => 268),
  (x => 353, y => 268),
  (x => 354, y => 268),
  (x => 355, y => 268),
  (x => 356, y => 268),
  (x => 357, y => 268),
  (x => 358, y => 268),
  (x => 359, y => 268),
  (x => 376, y => 268),
  (x => 377, y => 268),
  (x => 378, y => 268),
  (x => 265, y => 269),
  (x => 266, y => 269),
  (x => 267, y => 269),
  (x => 268, y => 269),
  (x => 274, y => 269),
  (x => 275, y => 269),
  (x => 276, y => 269),
  (x => 277, y => 269),
  (x => 278, y => 269),
  (x => 284, y => 269),
  (x => 285, y => 269),
  (x => 286, y => 269),
  (x => 287, y => 269),
  (x => 296, y => 269),
  (x => 297, y => 269),
  (x => 298, y => 269),
  (x => 306, y => 269),
  (x => 307, y => 269),
  (x => 312, y => 269),
  (x => 313, y => 269),
  (x => 314, y => 269),
  (x => 326, y => 269),
  (x => 327, y => 269),
  (x => 328, y => 269),
  (x => 350, y => 269),
  (x => 351, y => 269),
  (x => 352, y => 269),
  (x => 353, y => 269),
  (x => 354, y => 269),
  (x => 355, y => 269),
  (x => 356, y => 269),
  (x => 357, y => 269),
  (x => 358, y => 269),
  (x => 359, y => 269),
  (x => 376, y => 269),
  (x => 377, y => 269),
  (x => 378, y => 269),
  (x => 265, y => 270),
  (x => 266, y => 270),
  (x => 267, y => 270),
  (x => 268, y => 270),
  (x => 269, y => 270),
  (x => 270, y => 270),
  (x => 271, y => 270),
  (x => 272, y => 270),
  (x => 273, y => 270),
  (x => 274, y => 270),
  (x => 275, y => 270),
  (x => 276, y => 270),
  (x => 277, y => 270),
  (x => 284, y => 270),
  (x => 285, y => 270),
  (x => 286, y => 270),
  (x => 287, y => 270),
  (x => 296, y => 270),
  (x => 297, y => 270),
  (x => 298, y => 270),
  (x => 306, y => 270),
  (x => 307, y => 270),
  (x => 308, y => 270),
  (x => 312, y => 270),
  (x => 313, y => 270),
  (x => 314, y => 270),
  (x => 315, y => 270),
  (x => 326, y => 270),
  (x => 327, y => 270),
  (x => 328, y => 270),
  (x => 329, y => 270),
  (x => 350, y => 270),
  (x => 351, y => 270),
  (x => 352, y => 270),
  (x => 353, y => 270),
  (x => 354, y => 270),
  (x => 355, y => 270),
  (x => 356, y => 270),
  (x => 357, y => 270),
  (x => 358, y => 270),
  (x => 359, y => 270),
  (x => 360, y => 270),
  (x => 361, y => 270),
  (x => 362, y => 270),
  (x => 376, y => 270),
  (x => 377, y => 270),
  (x => 378, y => 270),
  (x => 265, y => 271),
  (x => 266, y => 271),
  (x => 267, y => 271),
  (x => 268, y => 271),
  (x => 269, y => 271),
  (x => 270, y => 271),
  (x => 271, y => 271),
  (x => 272, y => 271),
  (x => 273, y => 271),
  (x => 274, y => 271),
  (x => 275, y => 271),
  (x => 276, y => 271),
  (x => 284, y => 271),
  (x => 285, y => 271),
  (x => 286, y => 271),
  (x => 287, y => 271),
  (x => 296, y => 271),
  (x => 297, y => 271),
  (x => 298, y => 271),
  (x => 306, y => 271),
  (x => 307, y => 271),
  (x => 308, y => 271),
  (x => 312, y => 271),
  (x => 313, y => 271),
  (x => 314, y => 271),
  (x => 315, y => 271),
  (x => 316, y => 271),
  (x => 326, y => 271),
  (x => 327, y => 271),
  (x => 328, y => 271),
  (x => 329, y => 271),
  (x => 330, y => 271),
  (x => 350, y => 271),
  (x => 351, y => 271),
  (x => 352, y => 271),
  (x => 353, y => 271),
  (x => 358, y => 271),
  (x => 359, y => 271),
  (x => 360, y => 271),
  (x => 361, y => 271),
  (x => 362, y => 271),
  (x => 363, y => 271),
  (x => 376, y => 271),
  (x => 377, y => 271),
  (x => 378, y => 271),
  (x => 265, y => 272),
  (x => 266, y => 272),
  (x => 267, y => 272),
  (x => 268, y => 272),
  (x => 269, y => 272),
  (x => 270, y => 272),
  (x => 271, y => 272),
  (x => 272, y => 272),
  (x => 273, y => 272),
  (x => 274, y => 272),
  (x => 275, y => 272),
  (x => 284, y => 272),
  (x => 285, y => 272),
  (x => 286, y => 272),
  (x => 295, y => 272),
  (x => 296, y => 272),
  (x => 297, y => 272),
  (x => 298, y => 272),
  (x => 306, y => 272),
  (x => 307, y => 272),
  (x => 308, y => 272),
  (x => 313, y => 272),
  (x => 314, y => 272),
  (x => 315, y => 272),
  (x => 316, y => 272),
  (x => 317, y => 272),
  (x => 318, y => 272),
  (x => 327, y => 272),
  (x => 328, y => 272),
  (x => 329, y => 272),
  (x => 330, y => 272),
  (x => 331, y => 272),
  (x => 332, y => 272),
  (x => 350, y => 272),
  (x => 351, y => 272),
  (x => 352, y => 272),
  (x => 353, y => 272),
  (x => 360, y => 272),
  (x => 361, y => 272),
  (x => 362, y => 272),
  (x => 363, y => 272),
  (x => 364, y => 272),
  (x => 376, y => 272),
  (x => 377, y => 272),
  (x => 378, y => 272),
  (x => 265, y => 273),
  (x => 266, y => 273),
  (x => 267, y => 273),
  (x => 268, y => 273),
  (x => 269, y => 273),
  (x => 270, y => 273),
  (x => 271, y => 273),
  (x => 272, y => 273),
  (x => 273, y => 273),
  (x => 274, y => 273),
  (x => 284, y => 273),
  (x => 285, y => 273),
  (x => 286, y => 273),
  (x => 295, y => 273),
  (x => 296, y => 273),
  (x => 297, y => 273),
  (x => 298, y => 273),
  (x => 299, y => 273),
  (x => 300, y => 273),
  (x => 301, y => 273),
  (x => 302, y => 273),
  (x => 303, y => 273),
  (x => 304, y => 273),
  (x => 305, y => 273),
  (x => 306, y => 273),
  (x => 307, y => 273),
  (x => 308, y => 273),
  (x => 313, y => 273),
  (x => 314, y => 273),
  (x => 315, y => 273),
  (x => 316, y => 273),
  (x => 317, y => 273),
  (x => 318, y => 273),
  (x => 319, y => 273),
  (x => 320, y => 273),
  (x => 327, y => 273),
  (x => 328, y => 273),
  (x => 329, y => 273),
  (x => 330, y => 273),
  (x => 331, y => 273),
  (x => 332, y => 273),
  (x => 333, y => 273),
  (x => 350, y => 273),
  (x => 351, y => 273),
  (x => 352, y => 273),
  (x => 353, y => 273),
  (x => 361, y => 273),
  (x => 362, y => 273),
  (x => 363, y => 273),
  (x => 364, y => 273),
  (x => 376, y => 273),
  (x => 377, y => 273),
  (x => 378, y => 273),
  (x => 265, y => 274),
  (x => 266, y => 274),
  (x => 267, y => 274),
  (x => 268, y => 274),
  (x => 284, y => 274),
  (x => 285, y => 274),
  (x => 286, y => 274),
  (x => 295, y => 274),
  (x => 296, y => 274),
  (x => 297, y => 274),
  (x => 298, y => 274),
  (x => 299, y => 274),
  (x => 300, y => 274),
  (x => 301, y => 274),
  (x => 302, y => 274),
  (x => 303, y => 274),
  (x => 304, y => 274),
  (x => 305, y => 274),
  (x => 306, y => 274),
  (x => 307, y => 274),
  (x => 308, y => 274),
  (x => 314, y => 274),
  (x => 315, y => 274),
  (x => 316, y => 274),
  (x => 317, y => 274),
  (x => 318, y => 274),
  (x => 319, y => 274),
  (x => 320, y => 274),
  (x => 321, y => 274),
  (x => 328, y => 274),
  (x => 329, y => 274),
  (x => 330, y => 274),
  (x => 331, y => 274),
  (x => 332, y => 274),
  (x => 333, y => 274),
  (x => 334, y => 274),
  (x => 335, y => 274),
  (x => 350, y => 274),
  (x => 351, y => 274),
  (x => 352, y => 274),
  (x => 353, y => 274),
  (x => 361, y => 274),
  (x => 362, y => 274),
  (x => 363, y => 274),
  (x => 364, y => 274),
  (x => 376, y => 274),
  (x => 377, y => 274),
  (x => 378, y => 274),
  (x => 265, y => 275),
  (x => 266, y => 275),
  (x => 267, y => 275),
  (x => 268, y => 275),
  (x => 284, y => 275),
  (x => 285, y => 275),
  (x => 286, y => 275),
  (x => 295, y => 275),
  (x => 296, y => 275),
  (x => 297, y => 275),
  (x => 298, y => 275),
  (x => 300, y => 275),
  (x => 301, y => 275),
  (x => 302, y => 275),
  (x => 303, y => 275),
  (x => 304, y => 275),
  (x => 305, y => 275),
  (x => 306, y => 275),
  (x => 307, y => 275),
  (x => 308, y => 275),
  (x => 316, y => 275),
  (x => 317, y => 275),
  (x => 318, y => 275),
  (x => 319, y => 275),
  (x => 320, y => 275),
  (x => 321, y => 275),
  (x => 330, y => 275),
  (x => 331, y => 275),
  (x => 332, y => 275),
  (x => 333, y => 275),
  (x => 334, y => 275),
  (x => 335, y => 275),
  (x => 350, y => 275),
  (x => 351, y => 275),
  (x => 352, y => 275),
  (x => 353, y => 275),
  (x => 362, y => 275),
  (x => 363, y => 275),
  (x => 364, y => 275),
  (x => 376, y => 275),
  (x => 377, y => 275),
  (x => 378, y => 275),
  (x => 265, y => 276),
  (x => 266, y => 276),
  (x => 267, y => 276),
  (x => 268, y => 276),
  (x => 284, y => 276),
  (x => 285, y => 276),
  (x => 286, y => 276),
  (x => 295, y => 276),
  (x => 296, y => 276),
  (x => 297, y => 276),
  (x => 298, y => 276),
  (x => 318, y => 276),
  (x => 319, y => 276),
  (x => 320, y => 276),
  (x => 321, y => 276),
  (x => 322, y => 276),
  (x => 332, y => 276),
  (x => 333, y => 276),
  (x => 334, y => 276),
  (x => 335, y => 276),
  (x => 336, y => 276),
  (x => 350, y => 276),
  (x => 351, y => 276),
  (x => 352, y => 276),
  (x => 353, y => 276),
  (x => 362, y => 276),
  (x => 363, y => 276),
  (x => 364, y => 276),
  (x => 376, y => 276),
  (x => 377, y => 276),
  (x => 378, y => 276),
  (x => 265, y => 277),
  (x => 266, y => 277),
  (x => 267, y => 277),
  (x => 268, y => 277),
  (x => 284, y => 277),
  (x => 285, y => 277),
  (x => 286, y => 277),
  (x => 296, y => 277),
  (x => 297, y => 277),
  (x => 298, y => 277),
  (x => 319, y => 277),
  (x => 320, y => 277),
  (x => 321, y => 277),
  (x => 322, y => 277),
  (x => 333, y => 277),
  (x => 334, y => 277),
  (x => 335, y => 277),
  (x => 336, y => 277),
  (x => 350, y => 277),
  (x => 351, y => 277),
  (x => 352, y => 277),
  (x => 353, y => 277),
  (x => 361, y => 277),
  (x => 362, y => 277),
  (x => 363, y => 277),
  (x => 364, y => 277),
  (x => 376, y => 277),
  (x => 377, y => 277),
  (x => 378, y => 277),
  (x => 265, y => 278),
  (x => 266, y => 278),
  (x => 267, y => 278),
  (x => 268, y => 278),
  (x => 284, y => 278),
  (x => 285, y => 278),
  (x => 286, y => 278),
  (x => 296, y => 278),
  (x => 297, y => 278),
  (x => 298, y => 278),
  (x => 320, y => 278),
  (x => 321, y => 278),
  (x => 322, y => 278),
  (x => 334, y => 278),
  (x => 335, y => 278),
  (x => 336, y => 278),
  (x => 350, y => 278),
  (x => 351, y => 278),
  (x => 352, y => 278),
  (x => 353, y => 278),
  (x => 361, y => 278),
  (x => 362, y => 278),
  (x => 363, y => 278),
  (x => 364, y => 278),
  (x => 376, y => 278),
  (x => 377, y => 278),
  (x => 378, y => 278),
  (x => 265, y => 279),
  (x => 266, y => 279),
  (x => 267, y => 279),
  (x => 268, y => 279),
  (x => 284, y => 279),
  (x => 285, y => 279),
  (x => 286, y => 279),
  (x => 296, y => 279),
  (x => 297, y => 279),
  (x => 298, y => 279),
  (x => 299, y => 279),
  (x => 320, y => 279),
  (x => 321, y => 279),
  (x => 322, y => 279),
  (x => 333, y => 279),
  (x => 334, y => 279),
  (x => 335, y => 279),
  (x => 336, y => 279),
  (x => 350, y => 279),
  (x => 351, y => 279),
  (x => 352, y => 279),
  (x => 353, y => 279),
  (x => 360, y => 279),
  (x => 361, y => 279),
  (x => 362, y => 279),
  (x => 363, y => 279),
  (x => 364, y => 279),
  (x => 376, y => 279),
  (x => 377, y => 279),
  (x => 378, y => 279),
  (x => 265, y => 280),
  (x => 266, y => 280),
  (x => 267, y => 280),
  (x => 268, y => 280),
  (x => 284, y => 280),
  (x => 285, y => 280),
  (x => 286, y => 280),
  (x => 296, y => 280),
  (x => 297, y => 280),
  (x => 298, y => 280),
  (x => 299, y => 280),
  (x => 300, y => 280),
  (x => 307, y => 280),
  (x => 312, y => 280),
  (x => 319, y => 280),
  (x => 320, y => 280),
  (x => 321, y => 280),
  (x => 322, y => 280),
  (x => 326, y => 280),
  (x => 333, y => 280),
  (x => 334, y => 280),
  (x => 335, y => 280),
  (x => 350, y => 280),
  (x => 351, y => 280),
  (x => 352, y => 280),
  (x => 353, y => 280),
  (x => 354, y => 280),
  (x => 355, y => 280),
  (x => 356, y => 280),
  (x => 357, y => 280),
  (x => 358, y => 280),
  (x => 359, y => 280),
  (x => 360, y => 280),
  (x => 361, y => 280),
  (x => 362, y => 280),
  (x => 363, y => 280),
  (x => 376, y => 280),
  (x => 377, y => 280),
  (x => 378, y => 280),
  (x => 265, y => 281),
  (x => 266, y => 281),
  (x => 267, y => 281),
  (x => 268, y => 281),
  (x => 284, y => 281),
  (x => 285, y => 281),
  (x => 286, y => 281),
  (x => 297, y => 281),
  (x => 298, y => 281),
  (x => 299, y => 281),
  (x => 300, y => 281),
  (x => 301, y => 281),
  (x => 302, y => 281),
  (x => 303, y => 281),
  (x => 304, y => 281),
  (x => 305, y => 281),
  (x => 306, y => 281),
  (x => 307, y => 281),
  (x => 312, y => 281),
  (x => 313, y => 281),
  (x => 314, y => 281),
  (x => 315, y => 281),
  (x => 316, y => 281),
  (x => 317, y => 281),
  (x => 318, y => 281),
  (x => 319, y => 281),
  (x => 320, y => 281),
  (x => 321, y => 281),
  (x => 326, y => 281),
  (x => 327, y => 281),
  (x => 328, y => 281),
  (x => 329, y => 281),
  (x => 330, y => 281),
  (x => 331, y => 281),
  (x => 332, y => 281),
  (x => 333, y => 281),
  (x => 334, y => 281),
  (x => 335, y => 281),
  (x => 350, y => 281),
  (x => 351, y => 281),
  (x => 352, y => 281),
  (x => 353, y => 281),
  (x => 354, y => 281),
  (x => 355, y => 281),
  (x => 356, y => 281),
  (x => 357, y => 281),
  (x => 358, y => 281),
  (x => 359, y => 281),
  (x => 360, y => 281),
  (x => 361, y => 281),
  (x => 362, y => 281),
  (x => 363, y => 281),
  (x => 376, y => 281),
  (x => 377, y => 281),
  (x => 378, y => 281),
  (x => 265, y => 282),
  (x => 266, y => 282),
  (x => 267, y => 282),
  (x => 268, y => 282),
  (x => 284, y => 282),
  (x => 285, y => 282),
  (x => 286, y => 282),
  (x => 298, y => 282),
  (x => 299, y => 282),
  (x => 300, y => 282),
  (x => 301, y => 282),
  (x => 302, y => 282),
  (x => 303, y => 282),
  (x => 304, y => 282),
  (x => 305, y => 282),
  (x => 306, y => 282),
  (x => 307, y => 282),
  (x => 312, y => 282),
  (x => 313, y => 282),
  (x => 314, y => 282),
  (x => 315, y => 282),
  (x => 316, y => 282),
  (x => 317, y => 282),
  (x => 318, y => 282),
  (x => 319, y => 282),
  (x => 320, y => 282),
  (x => 326, y => 282),
  (x => 327, y => 282),
  (x => 328, y => 282),
  (x => 329, y => 282),
  (x => 330, y => 282),
  (x => 331, y => 282),
  (x => 332, y => 282),
  (x => 333, y => 282),
  (x => 334, y => 282),
  (x => 350, y => 282),
  (x => 351, y => 282),
  (x => 352, y => 282),
  (x => 353, y => 282),
  (x => 354, y => 282),
  (x => 355, y => 282),
  (x => 356, y => 282),
  (x => 357, y => 282),
  (x => 358, y => 282),
  (x => 359, y => 282),
  (x => 360, y => 282),
  (x => 361, y => 282),
  (x => 362, y => 282),
  (x => 376, y => 282),
  (x => 377, y => 282),
  (x => 378, y => 282),
  (x => 265, y => 283),
  (x => 266, y => 283),
  (x => 267, y => 283),
  (x => 268, y => 283),
  (x => 284, y => 283),
  (x => 285, y => 283),
  (x => 286, y => 283),
  (x => 299, y => 283),
  (x => 300, y => 283),
  (x => 301, y => 283),
  (x => 302, y => 283),
  (x => 303, y => 283),
  (x => 304, y => 283),
  (x => 305, y => 283),
  (x => 306, y => 283),
  (x => 312, y => 283),
  (x => 313, y => 283),
  (x => 314, y => 283),
  (x => 315, y => 283),
  (x => 316, y => 283),
  (x => 317, y => 283),
  (x => 318, y => 283),
  (x => 319, y => 283),
  (x => 326, y => 283),
  (x => 327, y => 283),
  (x => 328, y => 283),
  (x => 329, y => 283),
  (x => 330, y => 283),
  (x => 331, y => 283),
  (x => 332, y => 283),
  (x => 333, y => 283),
  (x => 350, y => 283),
  (x => 351, y => 283),
  (x => 352, y => 283),
  (x => 353, y => 283),
  (x => 354, y => 283),
  (x => 355, y => 283),
  (x => 356, y => 283),
  (x => 357, y => 283),
  (x => 358, y => 283),
  (x => 359, y => 283),
  (x => 360, y => 283),
  (x => 376, y => 283),
  (x => 377, y => 283),
  (x => 378, y => 283)
);
constant p1_end_screen: CoordPairArray(0 to 6548) := (
  (x => 177, y => 128),
  (x => 178, y => 128),
  (x => 179, y => 128),
  (x => 180, y => 128),
  (x => 181, y => 128),
  (x => 182, y => 128),
  (x => 183, y => 128),
  (x => 184, y => 128),
  (x => 185, y => 128),
  (x => 186, y => 128),
  (x => 187, y => 128),
  (x => 188, y => 128),
  (x => 337, y => 128),
  (x => 338, y => 128),
  (x => 339, y => 128),
  (x => 340, y => 128),
  (x => 341, y => 128),
  (x => 342, y => 128),
  (x => 343, y => 128),
  (x => 344, y => 128),
  (x => 345, y => 128),
  (x => 175, y => 129),
  (x => 176, y => 129),
  (x => 177, y => 129),
  (x => 178, y => 129),
  (x => 179, y => 129),
  (x => 180, y => 129),
  (x => 181, y => 129),
  (x => 182, y => 129),
  (x => 183, y => 129),
  (x => 184, y => 129),
  (x => 185, y => 129),
  (x => 186, y => 129),
  (x => 187, y => 129),
  (x => 188, y => 129),
  (x => 189, y => 129),
  (x => 190, y => 129),
  (x => 191, y => 129),
  (x => 334, y => 129),
  (x => 335, y => 129),
  (x => 336, y => 129),
  (x => 337, y => 129),
  (x => 338, y => 129),
  (x => 339, y => 129),
  (x => 340, y => 129),
  (x => 341, y => 129),
  (x => 342, y => 129),
  (x => 343, y => 129),
  (x => 344, y => 129),
  (x => 345, y => 129),
  (x => 346, y => 129),
  (x => 347, y => 129),
  (x => 173, y => 130),
  (x => 174, y => 130),
  (x => 175, y => 130),
  (x => 176, y => 130),
  (x => 177, y => 130),
  (x => 178, y => 130),
  (x => 179, y => 130),
  (x => 180, y => 130),
  (x => 181, y => 130),
  (x => 182, y => 130),
  (x => 183, y => 130),
  (x => 184, y => 130),
  (x => 185, y => 130),
  (x => 186, y => 130),
  (x => 187, y => 130),
  (x => 188, y => 130),
  (x => 189, y => 130),
  (x => 190, y => 130),
  (x => 191, y => 130),
  (x => 333, y => 130),
  (x => 334, y => 130),
  (x => 335, y => 130),
  (x => 336, y => 130),
  (x => 337, y => 130),
  (x => 338, y => 130),
  (x => 339, y => 130),
  (x => 340, y => 130),
  (x => 341, y => 130),
  (x => 342, y => 130),
  (x => 343, y => 130),
  (x => 344, y => 130),
  (x => 345, y => 130),
  (x => 346, y => 130),
  (x => 347, y => 130),
  (x => 348, y => 130),
  (x => 349, y => 130),
  (x => 171, y => 131),
  (x => 172, y => 131),
  (x => 173, y => 131),
  (x => 174, y => 131),
  (x => 175, y => 131),
  (x => 176, y => 131),
  (x => 177, y => 131),
  (x => 178, y => 131),
  (x => 179, y => 131),
  (x => 180, y => 131),
  (x => 181, y => 131),
  (x => 182, y => 131),
  (x => 183, y => 131),
  (x => 184, y => 131),
  (x => 185, y => 131),
  (x => 186, y => 131),
  (x => 187, y => 131),
  (x => 188, y => 131),
  (x => 189, y => 131),
  (x => 190, y => 131),
  (x => 191, y => 131),
  (x => 331, y => 131),
  (x => 332, y => 131),
  (x => 333, y => 131),
  (x => 334, y => 131),
  (x => 335, y => 131),
  (x => 336, y => 131),
  (x => 337, y => 131),
  (x => 338, y => 131),
  (x => 339, y => 131),
  (x => 340, y => 131),
  (x => 341, y => 131),
  (x => 342, y => 131),
  (x => 343, y => 131),
  (x => 344, y => 131),
  (x => 345, y => 131),
  (x => 346, y => 131),
  (x => 347, y => 131),
  (x => 348, y => 131),
  (x => 349, y => 131),
  (x => 350, y => 131),
  (x => 170, y => 132),
  (x => 171, y => 132),
  (x => 172, y => 132),
  (x => 173, y => 132),
  (x => 174, y => 132),
  (x => 175, y => 132),
  (x => 176, y => 132),
  (x => 177, y => 132),
  (x => 178, y => 132),
  (x => 179, y => 132),
  (x => 180, y => 132),
  (x => 181, y => 132),
  (x => 182, y => 132),
  (x => 183, y => 132),
  (x => 184, y => 132),
  (x => 185, y => 132),
  (x => 186, y => 132),
  (x => 187, y => 132),
  (x => 188, y => 132),
  (x => 189, y => 132),
  (x => 190, y => 132),
  (x => 191, y => 132),
  (x => 330, y => 132),
  (x => 331, y => 132),
  (x => 332, y => 132),
  (x => 333, y => 132),
  (x => 334, y => 132),
  (x => 335, y => 132),
  (x => 336, y => 132),
  (x => 337, y => 132),
  (x => 338, y => 132),
  (x => 339, y => 132),
  (x => 340, y => 132),
  (x => 341, y => 132),
  (x => 342, y => 132),
  (x => 343, y => 132),
  (x => 344, y => 132),
  (x => 345, y => 132),
  (x => 346, y => 132),
  (x => 347, y => 132),
  (x => 348, y => 132),
  (x => 349, y => 132),
  (x => 350, y => 132),
  (x => 351, y => 132),
  (x => 169, y => 133),
  (x => 170, y => 133),
  (x => 171, y => 133),
  (x => 172, y => 133),
  (x => 173, y => 133),
  (x => 174, y => 133),
  (x => 175, y => 133),
  (x => 176, y => 133),
  (x => 177, y => 133),
  (x => 178, y => 133),
  (x => 179, y => 133),
  (x => 180, y => 133),
  (x => 181, y => 133),
  (x => 182, y => 133),
  (x => 183, y => 133),
  (x => 184, y => 133),
  (x => 185, y => 133),
  (x => 186, y => 133),
  (x => 187, y => 133),
  (x => 188, y => 133),
  (x => 189, y => 133),
  (x => 190, y => 133),
  (x => 191, y => 133),
  (x => 329, y => 133),
  (x => 330, y => 133),
  (x => 331, y => 133),
  (x => 332, y => 133),
  (x => 333, y => 133),
  (x => 334, y => 133),
  (x => 335, y => 133),
  (x => 336, y => 133),
  (x => 337, y => 133),
  (x => 338, y => 133),
  (x => 339, y => 133),
  (x => 340, y => 133),
  (x => 341, y => 133),
  (x => 342, y => 133),
  (x => 343, y => 133),
  (x => 344, y => 133),
  (x => 345, y => 133),
  (x => 346, y => 133),
  (x => 347, y => 133),
  (x => 348, y => 133),
  (x => 349, y => 133),
  (x => 350, y => 133),
  (x => 351, y => 133),
  (x => 352, y => 133),
  (x => 168, y => 134),
  (x => 169, y => 134),
  (x => 170, y => 134),
  (x => 171, y => 134),
  (x => 172, y => 134),
  (x => 173, y => 134),
  (x => 174, y => 134),
  (x => 175, y => 134),
  (x => 176, y => 134),
  (x => 177, y => 134),
  (x => 178, y => 134),
  (x => 179, y => 134),
  (x => 180, y => 134),
  (x => 181, y => 134),
  (x => 182, y => 134),
  (x => 183, y => 134),
  (x => 184, y => 134),
  (x => 185, y => 134),
  (x => 186, y => 134),
  (x => 187, y => 134),
  (x => 188, y => 134),
  (x => 189, y => 134),
  (x => 190, y => 134),
  (x => 191, y => 134),
  (x => 329, y => 134),
  (x => 330, y => 134),
  (x => 331, y => 134),
  (x => 332, y => 134),
  (x => 333, y => 134),
  (x => 334, y => 134),
  (x => 335, y => 134),
  (x => 336, y => 134),
  (x => 337, y => 134),
  (x => 338, y => 134),
  (x => 339, y => 134),
  (x => 340, y => 134),
  (x => 341, y => 134),
  (x => 342, y => 134),
  (x => 343, y => 134),
  (x => 344, y => 134),
  (x => 345, y => 134),
  (x => 346, y => 134),
  (x => 347, y => 134),
  (x => 348, y => 134),
  (x => 349, y => 134),
  (x => 350, y => 134),
  (x => 351, y => 134),
  (x => 352, y => 134),
  (x => 353, y => 134),
  (x => 167, y => 135),
  (x => 168, y => 135),
  (x => 169, y => 135),
  (x => 170, y => 135),
  (x => 171, y => 135),
  (x => 172, y => 135),
  (x => 173, y => 135),
  (x => 174, y => 135),
  (x => 175, y => 135),
  (x => 176, y => 135),
  (x => 177, y => 135),
  (x => 178, y => 135),
  (x => 179, y => 135),
  (x => 180, y => 135),
  (x => 181, y => 135),
  (x => 182, y => 135),
  (x => 183, y => 135),
  (x => 184, y => 135),
  (x => 185, y => 135),
  (x => 186, y => 135),
  (x => 187, y => 135),
  (x => 188, y => 135),
  (x => 189, y => 135),
  (x => 190, y => 135),
  (x => 191, y => 135),
  (x => 328, y => 135),
  (x => 329, y => 135),
  (x => 330, y => 135),
  (x => 331, y => 135),
  (x => 332, y => 135),
  (x => 333, y => 135),
  (x => 334, y => 135),
  (x => 335, y => 135),
  (x => 336, y => 135),
  (x => 337, y => 135),
  (x => 338, y => 135),
  (x => 339, y => 135),
  (x => 340, y => 135),
  (x => 341, y => 135),
  (x => 342, y => 135),
  (x => 343, y => 135),
  (x => 344, y => 135),
  (x => 345, y => 135),
  (x => 346, y => 135),
  (x => 347, y => 135),
  (x => 348, y => 135),
  (x => 349, y => 135),
  (x => 350, y => 135),
  (x => 351, y => 135),
  (x => 352, y => 135),
  (x => 353, y => 135),
  (x => 354, y => 135),
  (x => 167, y => 136),
  (x => 168, y => 136),
  (x => 169, y => 136),
  (x => 170, y => 136),
  (x => 171, y => 136),
  (x => 172, y => 136),
  (x => 173, y => 136),
  (x => 174, y => 136),
  (x => 175, y => 136),
  (x => 176, y => 136),
  (x => 177, y => 136),
  (x => 178, y => 136),
  (x => 188, y => 136),
  (x => 189, y => 136),
  (x => 190, y => 136),
  (x => 191, y => 136),
  (x => 327, y => 136),
  (x => 328, y => 136),
  (x => 329, y => 136),
  (x => 330, y => 136),
  (x => 331, y => 136),
  (x => 332, y => 136),
  (x => 333, y => 136),
  (x => 334, y => 136),
  (x => 335, y => 136),
  (x => 336, y => 136),
  (x => 337, y => 136),
  (x => 338, y => 136),
  (x => 344, y => 136),
  (x => 345, y => 136),
  (x => 346, y => 136),
  (x => 347, y => 136),
  (x => 348, y => 136),
  (x => 349, y => 136),
  (x => 350, y => 136),
  (x => 351, y => 136),
  (x => 352, y => 136),
  (x => 353, y => 136),
  (x => 354, y => 136),
  (x => 166, y => 137),
  (x => 167, y => 137),
  (x => 168, y => 137),
  (x => 169, y => 137),
  (x => 170, y => 137),
  (x => 171, y => 137),
  (x => 172, y => 137),
  (x => 173, y => 137),
  (x => 174, y => 137),
  (x => 175, y => 137),
  (x => 176, y => 137),
  (x => 190, y => 137),
  (x => 191, y => 137),
  (x => 327, y => 137),
  (x => 328, y => 137),
  (x => 329, y => 137),
  (x => 330, y => 137),
  (x => 331, y => 137),
  (x => 332, y => 137),
  (x => 333, y => 137),
  (x => 334, y => 137),
  (x => 335, y => 137),
  (x => 336, y => 137),
  (x => 346, y => 137),
  (x => 347, y => 137),
  (x => 348, y => 137),
  (x => 349, y => 137),
  (x => 350, y => 137),
  (x => 351, y => 137),
  (x => 352, y => 137),
  (x => 353, y => 137),
  (x => 354, y => 137),
  (x => 355, y => 137),
  (x => 166, y => 138),
  (x => 167, y => 138),
  (x => 168, y => 138),
  (x => 169, y => 138),
  (x => 170, y => 138),
  (x => 171, y => 138),
  (x => 172, y => 138),
  (x => 173, y => 138),
  (x => 174, y => 138),
  (x => 326, y => 138),
  (x => 327, y => 138),
  (x => 328, y => 138),
  (x => 329, y => 138),
  (x => 330, y => 138),
  (x => 331, y => 138),
  (x => 332, y => 138),
  (x => 333, y => 138),
  (x => 334, y => 138),
  (x => 347, y => 138),
  (x => 348, y => 138),
  (x => 349, y => 138),
  (x => 350, y => 138),
  (x => 351, y => 138),
  (x => 352, y => 138),
  (x => 353, y => 138),
  (x => 354, y => 138),
  (x => 355, y => 138),
  (x => 165, y => 139),
  (x => 166, y => 139),
  (x => 167, y => 139),
  (x => 168, y => 139),
  (x => 169, y => 139),
  (x => 170, y => 139),
  (x => 171, y => 139),
  (x => 172, y => 139),
  (x => 173, y => 139),
  (x => 326, y => 139),
  (x => 327, y => 139),
  (x => 328, y => 139),
  (x => 329, y => 139),
  (x => 330, y => 139),
  (x => 331, y => 139),
  (x => 332, y => 139),
  (x => 333, y => 139),
  (x => 334, y => 139),
  (x => 348, y => 139),
  (x => 349, y => 139),
  (x => 350, y => 139),
  (x => 351, y => 139),
  (x => 352, y => 139),
  (x => 353, y => 139),
  (x => 354, y => 139),
  (x => 355, y => 139),
  (x => 356, y => 139),
  (x => 165, y => 140),
  (x => 166, y => 140),
  (x => 167, y => 140),
  (x => 168, y => 140),
  (x => 169, y => 140),
  (x => 170, y => 140),
  (x => 171, y => 140),
  (x => 172, y => 140),
  (x => 325, y => 140),
  (x => 326, y => 140),
  (x => 327, y => 140),
  (x => 328, y => 140),
  (x => 329, y => 140),
  (x => 330, y => 140),
  (x => 331, y => 140),
  (x => 332, y => 140),
  (x => 333, y => 140),
  (x => 348, y => 140),
  (x => 349, y => 140),
  (x => 350, y => 140),
  (x => 351, y => 140),
  (x => 352, y => 140),
  (x => 353, y => 140),
  (x => 354, y => 140),
  (x => 355, y => 140),
  (x => 356, y => 140),
  (x => 164, y => 141),
  (x => 165, y => 141),
  (x => 166, y => 141),
  (x => 167, y => 141),
  (x => 168, y => 141),
  (x => 169, y => 141),
  (x => 170, y => 141),
  (x => 171, y => 141),
  (x => 172, y => 141),
  (x => 325, y => 141),
  (x => 326, y => 141),
  (x => 327, y => 141),
  (x => 328, y => 141),
  (x => 329, y => 141),
  (x => 330, y => 141),
  (x => 331, y => 141),
  (x => 332, y => 141),
  (x => 349, y => 141),
  (x => 350, y => 141),
  (x => 351, y => 141),
  (x => 352, y => 141),
  (x => 353, y => 141),
  (x => 354, y => 141),
  (x => 355, y => 141),
  (x => 356, y => 141),
  (x => 164, y => 142),
  (x => 165, y => 142),
  (x => 166, y => 142),
  (x => 167, y => 142),
  (x => 168, y => 142),
  (x => 169, y => 142),
  (x => 170, y => 142),
  (x => 171, y => 142),
  (x => 210, y => 142),
  (x => 211, y => 142),
  (x => 212, y => 142),
  (x => 213, y => 142),
  (x => 214, y => 142),
  (x => 246, y => 142),
  (x => 247, y => 142),
  (x => 248, y => 142),
  (x => 263, y => 142),
  (x => 264, y => 142),
  (x => 265, y => 142),
  (x => 290, y => 142),
  (x => 291, y => 142),
  (x => 292, y => 142),
  (x => 293, y => 142),
  (x => 325, y => 142),
  (x => 326, y => 142),
  (x => 327, y => 142),
  (x => 328, y => 142),
  (x => 329, y => 142),
  (x => 330, y => 142),
  (x => 331, y => 142),
  (x => 332, y => 142),
  (x => 350, y => 142),
  (x => 351, y => 142),
  (x => 352, y => 142),
  (x => 353, y => 142),
  (x => 354, y => 142),
  (x => 355, y => 142),
  (x => 356, y => 142),
  (x => 357, y => 142),
  (x => 404, y => 142),
  (x => 405, y => 142),
  (x => 406, y => 142),
  (x => 407, y => 142),
  (x => 438, y => 142),
  (x => 439, y => 142),
  (x => 164, y => 143),
  (x => 165, y => 143),
  (x => 166, y => 143),
  (x => 167, y => 143),
  (x => 168, y => 143),
  (x => 169, y => 143),
  (x => 170, y => 143),
  (x => 171, y => 143),
  (x => 206, y => 143),
  (x => 207, y => 143),
  (x => 208, y => 143),
  (x => 209, y => 143),
  (x => 210, y => 143),
  (x => 211, y => 143),
  (x => 212, y => 143),
  (x => 213, y => 143),
  (x => 214, y => 143),
  (x => 215, y => 143),
  (x => 216, y => 143),
  (x => 217, y => 143),
  (x => 231, y => 143),
  (x => 232, y => 143),
  (x => 233, y => 143),
  (x => 234, y => 143),
  (x => 235, y => 143),
  (x => 236, y => 143),
  (x => 237, y => 143),
  (x => 243, y => 143),
  (x => 244, y => 143),
  (x => 245, y => 143),
  (x => 246, y => 143),
  (x => 247, y => 143),
  (x => 248, y => 143),
  (x => 249, y => 143),
  (x => 250, y => 143),
  (x => 251, y => 143),
  (x => 260, y => 143),
  (x => 261, y => 143),
  (x => 262, y => 143),
  (x => 263, y => 143),
  (x => 264, y => 143),
  (x => 265, y => 143),
  (x => 266, y => 143),
  (x => 267, y => 143),
  (x => 268, y => 143),
  (x => 287, y => 143),
  (x => 288, y => 143),
  (x => 289, y => 143),
  (x => 290, y => 143),
  (x => 291, y => 143),
  (x => 292, y => 143),
  (x => 293, y => 143),
  (x => 294, y => 143),
  (x => 295, y => 143),
  (x => 296, y => 143),
  (x => 324, y => 143),
  (x => 325, y => 143),
  (x => 326, y => 143),
  (x => 327, y => 143),
  (x => 328, y => 143),
  (x => 329, y => 143),
  (x => 330, y => 143),
  (x => 331, y => 143),
  (x => 350, y => 143),
  (x => 351, y => 143),
  (x => 352, y => 143),
  (x => 353, y => 143),
  (x => 354, y => 143),
  (x => 355, y => 143),
  (x => 356, y => 143),
  (x => 357, y => 143),
  (x => 362, y => 143),
  (x => 363, y => 143),
  (x => 364, y => 143),
  (x => 365, y => 143),
  (x => 366, y => 143),
  (x => 367, y => 143),
  (x => 368, y => 143),
  (x => 369, y => 143),
  (x => 382, y => 143),
  (x => 383, y => 143),
  (x => 384, y => 143),
  (x => 385, y => 143),
  (x => 386, y => 143),
  (x => 387, y => 143),
  (x => 388, y => 143),
  (x => 389, y => 143),
  (x => 401, y => 143),
  (x => 402, y => 143),
  (x => 403, y => 143),
  (x => 404, y => 143),
  (x => 405, y => 143),
  (x => 406, y => 143),
  (x => 407, y => 143),
  (x => 408, y => 143),
  (x => 409, y => 143),
  (x => 410, y => 143),
  (x => 424, y => 143),
  (x => 425, y => 143),
  (x => 426, y => 143),
  (x => 427, y => 143),
  (x => 428, y => 143),
  (x => 429, y => 143),
  (x => 430, y => 143),
  (x => 436, y => 143),
  (x => 437, y => 143),
  (x => 438, y => 143),
  (x => 439, y => 143),
  (x => 163, y => 144),
  (x => 164, y => 144),
  (x => 165, y => 144),
  (x => 166, y => 144),
  (x => 167, y => 144),
  (x => 168, y => 144),
  (x => 169, y => 144),
  (x => 170, y => 144),
  (x => 204, y => 144),
  (x => 205, y => 144),
  (x => 206, y => 144),
  (x => 207, y => 144),
  (x => 208, y => 144),
  (x => 209, y => 144),
  (x => 210, y => 144),
  (x => 211, y => 144),
  (x => 212, y => 144),
  (x => 213, y => 144),
  (x => 214, y => 144),
  (x => 215, y => 144),
  (x => 216, y => 144),
  (x => 217, y => 144),
  (x => 218, y => 144),
  (x => 231, y => 144),
  (x => 232, y => 144),
  (x => 233, y => 144),
  (x => 234, y => 144),
  (x => 235, y => 144),
  (x => 236, y => 144),
  (x => 237, y => 144),
  (x => 242, y => 144),
  (x => 243, y => 144),
  (x => 244, y => 144),
  (x => 245, y => 144),
  (x => 246, y => 144),
  (x => 247, y => 144),
  (x => 248, y => 144),
  (x => 249, y => 144),
  (x => 250, y => 144),
  (x => 251, y => 144),
  (x => 252, y => 144),
  (x => 259, y => 144),
  (x => 260, y => 144),
  (x => 261, y => 144),
  (x => 262, y => 144),
  (x => 263, y => 144),
  (x => 264, y => 144),
  (x => 265, y => 144),
  (x => 266, y => 144),
  (x => 267, y => 144),
  (x => 268, y => 144),
  (x => 269, y => 144),
  (x => 285, y => 144),
  (x => 286, y => 144),
  (x => 287, y => 144),
  (x => 288, y => 144),
  (x => 289, y => 144),
  (x => 290, y => 144),
  (x => 291, y => 144),
  (x => 292, y => 144),
  (x => 293, y => 144),
  (x => 294, y => 144),
  (x => 295, y => 144),
  (x => 296, y => 144),
  (x => 297, y => 144),
  (x => 324, y => 144),
  (x => 325, y => 144),
  (x => 326, y => 144),
  (x => 327, y => 144),
  (x => 328, y => 144),
  (x => 329, y => 144),
  (x => 330, y => 144),
  (x => 331, y => 144),
  (x => 350, y => 144),
  (x => 351, y => 144),
  (x => 352, y => 144),
  (x => 353, y => 144),
  (x => 354, y => 144),
  (x => 355, y => 144),
  (x => 356, y => 144),
  (x => 357, y => 144),
  (x => 363, y => 144),
  (x => 364, y => 144),
  (x => 365, y => 144),
  (x => 366, y => 144),
  (x => 367, y => 144),
  (x => 368, y => 144),
  (x => 369, y => 144),
  (x => 382, y => 144),
  (x => 383, y => 144),
  (x => 384, y => 144),
  (x => 385, y => 144),
  (x => 386, y => 144),
  (x => 387, y => 144),
  (x => 388, y => 144),
  (x => 400, y => 144),
  (x => 401, y => 144),
  (x => 402, y => 144),
  (x => 403, y => 144),
  (x => 404, y => 144),
  (x => 405, y => 144),
  (x => 406, y => 144),
  (x => 407, y => 144),
  (x => 408, y => 144),
  (x => 409, y => 144),
  (x => 410, y => 144),
  (x => 411, y => 144),
  (x => 412, y => 144),
  (x => 424, y => 144),
  (x => 425, y => 144),
  (x => 426, y => 144),
  (x => 427, y => 144),
  (x => 428, y => 144),
  (x => 429, y => 144),
  (x => 430, y => 144),
  (x => 435, y => 144),
  (x => 436, y => 144),
  (x => 437, y => 144),
  (x => 438, y => 144),
  (x => 439, y => 144),
  (x => 163, y => 145),
  (x => 164, y => 145),
  (x => 165, y => 145),
  (x => 166, y => 145),
  (x => 167, y => 145),
  (x => 168, y => 145),
  (x => 169, y => 145),
  (x => 170, y => 145),
  (x => 203, y => 145),
  (x => 204, y => 145),
  (x => 205, y => 145),
  (x => 206, y => 145),
  (x => 207, y => 145),
  (x => 208, y => 145),
  (x => 209, y => 145),
  (x => 210, y => 145),
  (x => 211, y => 145),
  (x => 212, y => 145),
  (x => 213, y => 145),
  (x => 214, y => 145),
  (x => 215, y => 145),
  (x => 216, y => 145),
  (x => 217, y => 145),
  (x => 218, y => 145),
  (x => 219, y => 145),
  (x => 231, y => 145),
  (x => 232, y => 145),
  (x => 233, y => 145),
  (x => 234, y => 145),
  (x => 235, y => 145),
  (x => 236, y => 145),
  (x => 237, y => 145),
  (x => 241, y => 145),
  (x => 242, y => 145),
  (x => 243, y => 145),
  (x => 244, y => 145),
  (x => 245, y => 145),
  (x => 246, y => 145),
  (x => 247, y => 145),
  (x => 248, y => 145),
  (x => 249, y => 145),
  (x => 250, y => 145),
  (x => 251, y => 145),
  (x => 252, y => 145),
  (x => 258, y => 145),
  (x => 259, y => 145),
  (x => 260, y => 145),
  (x => 261, y => 145),
  (x => 262, y => 145),
  (x => 263, y => 145),
  (x => 264, y => 145),
  (x => 265, y => 145),
  (x => 266, y => 145),
  (x => 267, y => 145),
  (x => 268, y => 145),
  (x => 269, y => 145),
  (x => 284, y => 145),
  (x => 285, y => 145),
  (x => 286, y => 145),
  (x => 287, y => 145),
  (x => 288, y => 145),
  (x => 289, y => 145),
  (x => 290, y => 145),
  (x => 291, y => 145),
  (x => 292, y => 145),
  (x => 293, y => 145),
  (x => 294, y => 145),
  (x => 295, y => 145),
  (x => 296, y => 145),
  (x => 297, y => 145),
  (x => 298, y => 145),
  (x => 324, y => 145),
  (x => 325, y => 145),
  (x => 326, y => 145),
  (x => 327, y => 145),
  (x => 328, y => 145),
  (x => 329, y => 145),
  (x => 330, y => 145),
  (x => 331, y => 145),
  (x => 350, y => 145),
  (x => 351, y => 145),
  (x => 352, y => 145),
  (x => 353, y => 145),
  (x => 354, y => 145),
  (x => 355, y => 145),
  (x => 356, y => 145),
  (x => 357, y => 145),
  (x => 363, y => 145),
  (x => 364, y => 145),
  (x => 365, y => 145),
  (x => 366, y => 145),
  (x => 367, y => 145),
  (x => 368, y => 145),
  (x => 369, y => 145),
  (x => 382, y => 145),
  (x => 383, y => 145),
  (x => 384, y => 145),
  (x => 385, y => 145),
  (x => 386, y => 145),
  (x => 387, y => 145),
  (x => 388, y => 145),
  (x => 399, y => 145),
  (x => 400, y => 145),
  (x => 401, y => 145),
  (x => 402, y => 145),
  (x => 403, y => 145),
  (x => 404, y => 145),
  (x => 405, y => 145),
  (x => 406, y => 145),
  (x => 407, y => 145),
  (x => 408, y => 145),
  (x => 409, y => 145),
  (x => 410, y => 145),
  (x => 411, y => 145),
  (x => 412, y => 145),
  (x => 413, y => 145),
  (x => 424, y => 145),
  (x => 425, y => 145),
  (x => 426, y => 145),
  (x => 427, y => 145),
  (x => 428, y => 145),
  (x => 429, y => 145),
  (x => 430, y => 145),
  (x => 434, y => 145),
  (x => 435, y => 145),
  (x => 436, y => 145),
  (x => 437, y => 145),
  (x => 438, y => 145),
  (x => 439, y => 145),
  (x => 163, y => 146),
  (x => 164, y => 146),
  (x => 165, y => 146),
  (x => 166, y => 146),
  (x => 167, y => 146),
  (x => 168, y => 146),
  (x => 169, y => 146),
  (x => 170, y => 146),
  (x => 203, y => 146),
  (x => 204, y => 146),
  (x => 205, y => 146),
  (x => 206, y => 146),
  (x => 207, y => 146),
  (x => 208, y => 146),
  (x => 209, y => 146),
  (x => 210, y => 146),
  (x => 211, y => 146),
  (x => 212, y => 146),
  (x => 213, y => 146),
  (x => 214, y => 146),
  (x => 215, y => 146),
  (x => 216, y => 146),
  (x => 217, y => 146),
  (x => 218, y => 146),
  (x => 219, y => 146),
  (x => 220, y => 146),
  (x => 231, y => 146),
  (x => 232, y => 146),
  (x => 233, y => 146),
  (x => 234, y => 146),
  (x => 235, y => 146),
  (x => 236, y => 146),
  (x => 237, y => 146),
  (x => 240, y => 146),
  (x => 241, y => 146),
  (x => 242, y => 146),
  (x => 243, y => 146),
  (x => 244, y => 146),
  (x => 245, y => 146),
  (x => 246, y => 146),
  (x => 247, y => 146),
  (x => 248, y => 146),
  (x => 249, y => 146),
  (x => 250, y => 146),
  (x => 251, y => 146),
  (x => 252, y => 146),
  (x => 253, y => 146),
  (x => 257, y => 146),
  (x => 258, y => 146),
  (x => 259, y => 146),
  (x => 260, y => 146),
  (x => 261, y => 146),
  (x => 262, y => 146),
  (x => 263, y => 146),
  (x => 264, y => 146),
  (x => 265, y => 146),
  (x => 266, y => 146),
  (x => 267, y => 146),
  (x => 268, y => 146),
  (x => 269, y => 146),
  (x => 270, y => 146),
  (x => 283, y => 146),
  (x => 284, y => 146),
  (x => 285, y => 146),
  (x => 286, y => 146),
  (x => 287, y => 146),
  (x => 288, y => 146),
  (x => 289, y => 146),
  (x => 290, y => 146),
  (x => 291, y => 146),
  (x => 292, y => 146),
  (x => 293, y => 146),
  (x => 294, y => 146),
  (x => 295, y => 146),
  (x => 296, y => 146),
  (x => 297, y => 146),
  (x => 298, y => 146),
  (x => 299, y => 146),
  (x => 324, y => 146),
  (x => 325, y => 146),
  (x => 326, y => 146),
  (x => 327, y => 146),
  (x => 328, y => 146),
  (x => 329, y => 146),
  (x => 330, y => 146),
  (x => 351, y => 146),
  (x => 352, y => 146),
  (x => 353, y => 146),
  (x => 354, y => 146),
  (x => 355, y => 146),
  (x => 356, y => 146),
  (x => 357, y => 146),
  (x => 363, y => 146),
  (x => 364, y => 146),
  (x => 365, y => 146),
  (x => 366, y => 146),
  (x => 367, y => 146),
  (x => 368, y => 146),
  (x => 369, y => 146),
  (x => 370, y => 146),
  (x => 382, y => 146),
  (x => 383, y => 146),
  (x => 384, y => 146),
  (x => 385, y => 146),
  (x => 386, y => 146),
  (x => 387, y => 146),
  (x => 388, y => 146),
  (x => 398, y => 146),
  (x => 399, y => 146),
  (x => 400, y => 146),
  (x => 401, y => 146),
  (x => 402, y => 146),
  (x => 403, y => 146),
  (x => 404, y => 146),
  (x => 405, y => 146),
  (x => 406, y => 146),
  (x => 407, y => 146),
  (x => 408, y => 146),
  (x => 409, y => 146),
  (x => 410, y => 146),
  (x => 411, y => 146),
  (x => 412, y => 146),
  (x => 413, y => 146),
  (x => 414, y => 146),
  (x => 424, y => 146),
  (x => 425, y => 146),
  (x => 426, y => 146),
  (x => 427, y => 146),
  (x => 428, y => 146),
  (x => 429, y => 146),
  (x => 430, y => 146),
  (x => 434, y => 146),
  (x => 435, y => 146),
  (x => 436, y => 146),
  (x => 437, y => 146),
  (x => 438, y => 146),
  (x => 439, y => 146),
  (x => 163, y => 147),
  (x => 164, y => 147),
  (x => 165, y => 147),
  (x => 166, y => 147),
  (x => 167, y => 147),
  (x => 168, y => 147),
  (x => 169, y => 147),
  (x => 203, y => 147),
  (x => 204, y => 147),
  (x => 205, y => 147),
  (x => 206, y => 147),
  (x => 207, y => 147),
  (x => 208, y => 147),
  (x => 209, y => 147),
  (x => 210, y => 147),
  (x => 211, y => 147),
  (x => 212, y => 147),
  (x => 213, y => 147),
  (x => 214, y => 147),
  (x => 215, y => 147),
  (x => 216, y => 147),
  (x => 217, y => 147),
  (x => 218, y => 147),
  (x => 219, y => 147),
  (x => 220, y => 147),
  (x => 231, y => 147),
  (x => 232, y => 147),
  (x => 233, y => 147),
  (x => 234, y => 147),
  (x => 235, y => 147),
  (x => 236, y => 147),
  (x => 237, y => 147),
  (x => 240, y => 147),
  (x => 241, y => 147),
  (x => 242, y => 147),
  (x => 243, y => 147),
  (x => 244, y => 147),
  (x => 245, y => 147),
  (x => 246, y => 147),
  (x => 247, y => 147),
  (x => 248, y => 147),
  (x => 249, y => 147),
  (x => 250, y => 147),
  (x => 251, y => 147),
  (x => 252, y => 147),
  (x => 253, y => 147),
  (x => 257, y => 147),
  (x => 258, y => 147),
  (x => 259, y => 147),
  (x => 260, y => 147),
  (x => 261, y => 147),
  (x => 262, y => 147),
  (x => 263, y => 147),
  (x => 264, y => 147),
  (x => 265, y => 147),
  (x => 266, y => 147),
  (x => 267, y => 147),
  (x => 268, y => 147),
  (x => 269, y => 147),
  (x => 270, y => 147),
  (x => 282, y => 147),
  (x => 283, y => 147),
  (x => 284, y => 147),
  (x => 285, y => 147),
  (x => 286, y => 147),
  (x => 287, y => 147),
  (x => 288, y => 147),
  (x => 289, y => 147),
  (x => 290, y => 147),
  (x => 291, y => 147),
  (x => 292, y => 147),
  (x => 293, y => 147),
  (x => 294, y => 147),
  (x => 295, y => 147),
  (x => 296, y => 147),
  (x => 297, y => 147),
  (x => 298, y => 147),
  (x => 299, y => 147),
  (x => 300, y => 147),
  (x => 324, y => 147),
  (x => 325, y => 147),
  (x => 326, y => 147),
  (x => 327, y => 147),
  (x => 328, y => 147),
  (x => 329, y => 147),
  (x => 330, y => 147),
  (x => 351, y => 147),
  (x => 352, y => 147),
  (x => 353, y => 147),
  (x => 354, y => 147),
  (x => 355, y => 147),
  (x => 356, y => 147),
  (x => 357, y => 147),
  (x => 358, y => 147),
  (x => 364, y => 147),
  (x => 365, y => 147),
  (x => 366, y => 147),
  (x => 367, y => 147),
  (x => 368, y => 147),
  (x => 369, y => 147),
  (x => 370, y => 147),
  (x => 382, y => 147),
  (x => 383, y => 147),
  (x => 384, y => 147),
  (x => 385, y => 147),
  (x => 386, y => 147),
  (x => 387, y => 147),
  (x => 388, y => 147),
  (x => 397, y => 147),
  (x => 398, y => 147),
  (x => 399, y => 147),
  (x => 400, y => 147),
  (x => 401, y => 147),
  (x => 402, y => 147),
  (x => 403, y => 147),
  (x => 404, y => 147),
  (x => 405, y => 147),
  (x => 406, y => 147),
  (x => 407, y => 147),
  (x => 408, y => 147),
  (x => 409, y => 147),
  (x => 410, y => 147),
  (x => 411, y => 147),
  (x => 412, y => 147),
  (x => 413, y => 147),
  (x => 414, y => 147),
  (x => 424, y => 147),
  (x => 425, y => 147),
  (x => 426, y => 147),
  (x => 427, y => 147),
  (x => 428, y => 147),
  (x => 429, y => 147),
  (x => 430, y => 147),
  (x => 433, y => 147),
  (x => 434, y => 147),
  (x => 435, y => 147),
  (x => 436, y => 147),
  (x => 437, y => 147),
  (x => 438, y => 147),
  (x => 439, y => 147),
  (x => 163, y => 148),
  (x => 164, y => 148),
  (x => 165, y => 148),
  (x => 166, y => 148),
  (x => 167, y => 148),
  (x => 168, y => 148),
  (x => 169, y => 148),
  (x => 203, y => 148),
  (x => 204, y => 148),
  (x => 205, y => 148),
  (x => 206, y => 148),
  (x => 207, y => 148),
  (x => 208, y => 148),
  (x => 213, y => 148),
  (x => 214, y => 148),
  (x => 215, y => 148),
  (x => 216, y => 148),
  (x => 217, y => 148),
  (x => 218, y => 148),
  (x => 219, y => 148),
  (x => 220, y => 148),
  (x => 221, y => 148),
  (x => 231, y => 148),
  (x => 232, y => 148),
  (x => 233, y => 148),
  (x => 234, y => 148),
  (x => 235, y => 148),
  (x => 236, y => 148),
  (x => 237, y => 148),
  (x => 239, y => 148),
  (x => 240, y => 148),
  (x => 241, y => 148),
  (x => 242, y => 148),
  (x => 243, y => 148),
  (x => 244, y => 148),
  (x => 245, y => 148),
  (x => 246, y => 148),
  (x => 247, y => 148),
  (x => 248, y => 148),
  (x => 249, y => 148),
  (x => 250, y => 148),
  (x => 251, y => 148),
  (x => 252, y => 148),
  (x => 253, y => 148),
  (x => 254, y => 148),
  (x => 256, y => 148),
  (x => 257, y => 148),
  (x => 258, y => 148),
  (x => 259, y => 148),
  (x => 260, y => 148),
  (x => 261, y => 148),
  (x => 262, y => 148),
  (x => 263, y => 148),
  (x => 264, y => 148),
  (x => 265, y => 148),
  (x => 266, y => 148),
  (x => 267, y => 148),
  (x => 268, y => 148),
  (x => 269, y => 148),
  (x => 270, y => 148),
  (x => 271, y => 148),
  (x => 282, y => 148),
  (x => 283, y => 148),
  (x => 284, y => 148),
  (x => 285, y => 148),
  (x => 286, y => 148),
  (x => 287, y => 148),
  (x => 288, y => 148),
  (x => 289, y => 148),
  (x => 293, y => 148),
  (x => 294, y => 148),
  (x => 295, y => 148),
  (x => 296, y => 148),
  (x => 297, y => 148),
  (x => 298, y => 148),
  (x => 299, y => 148),
  (x => 300, y => 148),
  (x => 324, y => 148),
  (x => 325, y => 148),
  (x => 326, y => 148),
  (x => 327, y => 148),
  (x => 328, y => 148),
  (x => 329, y => 148),
  (x => 330, y => 148),
  (x => 351, y => 148),
  (x => 352, y => 148),
  (x => 353, y => 148),
  (x => 354, y => 148),
  (x => 355, y => 148),
  (x => 356, y => 148),
  (x => 357, y => 148),
  (x => 358, y => 148),
  (x => 364, y => 148),
  (x => 365, y => 148),
  (x => 366, y => 148),
  (x => 367, y => 148),
  (x => 368, y => 148),
  (x => 369, y => 148),
  (x => 370, y => 148),
  (x => 382, y => 148),
  (x => 383, y => 148),
  (x => 384, y => 148),
  (x => 385, y => 148),
  (x => 386, y => 148),
  (x => 387, y => 148),
  (x => 396, y => 148),
  (x => 397, y => 148),
  (x => 398, y => 148),
  (x => 399, y => 148),
  (x => 400, y => 148),
  (x => 401, y => 148),
  (x => 402, y => 148),
  (x => 403, y => 148),
  (x => 404, y => 148),
  (x => 408, y => 148),
  (x => 409, y => 148),
  (x => 410, y => 148),
  (x => 411, y => 148),
  (x => 412, y => 148),
  (x => 413, y => 148),
  (x => 414, y => 148),
  (x => 415, y => 148),
  (x => 424, y => 148),
  (x => 425, y => 148),
  (x => 426, y => 148),
  (x => 427, y => 148),
  (x => 428, y => 148),
  (x => 429, y => 148),
  (x => 430, y => 148),
  (x => 433, y => 148),
  (x => 434, y => 148),
  (x => 435, y => 148),
  (x => 436, y => 148),
  (x => 437, y => 148),
  (x => 438, y => 148),
  (x => 439, y => 148),
  (x => 162, y => 149),
  (x => 163, y => 149),
  (x => 164, y => 149),
  (x => 165, y => 149),
  (x => 166, y => 149),
  (x => 167, y => 149),
  (x => 168, y => 149),
  (x => 169, y => 149),
  (x => 203, y => 149),
  (x => 204, y => 149),
  (x => 205, y => 149),
  (x => 215, y => 149),
  (x => 216, y => 149),
  (x => 217, y => 149),
  (x => 218, y => 149),
  (x => 219, y => 149),
  (x => 220, y => 149),
  (x => 221, y => 149),
  (x => 231, y => 149),
  (x => 232, y => 149),
  (x => 233, y => 149),
  (x => 234, y => 149),
  (x => 235, y => 149),
  (x => 236, y => 149),
  (x => 237, y => 149),
  (x => 238, y => 149),
  (x => 239, y => 149),
  (x => 240, y => 149),
  (x => 241, y => 149),
  (x => 245, y => 149),
  (x => 246, y => 149),
  (x => 247, y => 149),
  (x => 248, y => 149),
  (x => 249, y => 149),
  (x => 250, y => 149),
  (x => 251, y => 149),
  (x => 252, y => 149),
  (x => 253, y => 149),
  (x => 254, y => 149),
  (x => 255, y => 149),
  (x => 256, y => 149),
  (x => 257, y => 149),
  (x => 258, y => 149),
  (x => 262, y => 149),
  (x => 263, y => 149),
  (x => 264, y => 149),
  (x => 265, y => 149),
  (x => 266, y => 149),
  (x => 267, y => 149),
  (x => 268, y => 149),
  (x => 269, y => 149),
  (x => 270, y => 149),
  (x => 271, y => 149),
  (x => 281, y => 149),
  (x => 282, y => 149),
  (x => 283, y => 149),
  (x => 284, y => 149),
  (x => 285, y => 149),
  (x => 286, y => 149),
  (x => 287, y => 149),
  (x => 288, y => 149),
  (x => 295, y => 149),
  (x => 296, y => 149),
  (x => 297, y => 149),
  (x => 298, y => 149),
  (x => 299, y => 149),
  (x => 300, y => 149),
  (x => 301, y => 149),
  (x => 323, y => 149),
  (x => 324, y => 149),
  (x => 325, y => 149),
  (x => 326, y => 149),
  (x => 327, y => 149),
  (x => 328, y => 149),
  (x => 329, y => 149),
  (x => 330, y => 149),
  (x => 351, y => 149),
  (x => 352, y => 149),
  (x => 353, y => 149),
  (x => 354, y => 149),
  (x => 355, y => 149),
  (x => 356, y => 149),
  (x => 357, y => 149),
  (x => 358, y => 149),
  (x => 364, y => 149),
  (x => 365, y => 149),
  (x => 366, y => 149),
  (x => 367, y => 149),
  (x => 368, y => 149),
  (x => 369, y => 149),
  (x => 370, y => 149),
  (x => 381, y => 149),
  (x => 382, y => 149),
  (x => 383, y => 149),
  (x => 384, y => 149),
  (x => 385, y => 149),
  (x => 386, y => 149),
  (x => 387, y => 149),
  (x => 396, y => 149),
  (x => 397, y => 149),
  (x => 398, y => 149),
  (x => 399, y => 149),
  (x => 400, y => 149),
  (x => 401, y => 149),
  (x => 402, y => 149),
  (x => 409, y => 149),
  (x => 410, y => 149),
  (x => 411, y => 149),
  (x => 412, y => 149),
  (x => 413, y => 149),
  (x => 414, y => 149),
  (x => 415, y => 149),
  (x => 424, y => 149),
  (x => 425, y => 149),
  (x => 426, y => 149),
  (x => 427, y => 149),
  (x => 428, y => 149),
  (x => 429, y => 149),
  (x => 430, y => 149),
  (x => 431, y => 149),
  (x => 432, y => 149),
  (x => 433, y => 149),
  (x => 434, y => 149),
  (x => 435, y => 149),
  (x => 436, y => 149),
  (x => 437, y => 149),
  (x => 438, y => 149),
  (x => 439, y => 149),
  (x => 162, y => 150),
  (x => 163, y => 150),
  (x => 164, y => 150),
  (x => 165, y => 150),
  (x => 166, y => 150),
  (x => 167, y => 150),
  (x => 168, y => 150),
  (x => 169, y => 150),
  (x => 179, y => 150),
  (x => 180, y => 150),
  (x => 181, y => 150),
  (x => 182, y => 150),
  (x => 183, y => 150),
  (x => 184, y => 150),
  (x => 185, y => 150),
  (x => 186, y => 150),
  (x => 187, y => 150),
  (x => 188, y => 150),
  (x => 189, y => 150),
  (x => 190, y => 150),
  (x => 191, y => 150),
  (x => 192, y => 150),
  (x => 193, y => 150),
  (x => 203, y => 150),
  (x => 216, y => 150),
  (x => 217, y => 150),
  (x => 218, y => 150),
  (x => 219, y => 150),
  (x => 220, y => 150),
  (x => 221, y => 150),
  (x => 231, y => 150),
  (x => 232, y => 150),
  (x => 233, y => 150),
  (x => 234, y => 150),
  (x => 235, y => 150),
  (x => 236, y => 150),
  (x => 237, y => 150),
  (x => 238, y => 150),
  (x => 239, y => 150),
  (x => 246, y => 150),
  (x => 247, y => 150),
  (x => 248, y => 150),
  (x => 249, y => 150),
  (x => 250, y => 150),
  (x => 251, y => 150),
  (x => 252, y => 150),
  (x => 253, y => 150),
  (x => 254, y => 150),
  (x => 255, y => 150),
  (x => 256, y => 150),
  (x => 257, y => 150),
  (x => 264, y => 150),
  (x => 265, y => 150),
  (x => 266, y => 150),
  (x => 267, y => 150),
  (x => 268, y => 150),
  (x => 269, y => 150),
  (x => 270, y => 150),
  (x => 271, y => 150),
  (x => 281, y => 150),
  (x => 282, y => 150),
  (x => 283, y => 150),
  (x => 284, y => 150),
  (x => 285, y => 150),
  (x => 286, y => 150),
  (x => 287, y => 150),
  (x => 296, y => 150),
  (x => 297, y => 150),
  (x => 298, y => 150),
  (x => 299, y => 150),
  (x => 300, y => 150),
  (x => 301, y => 150),
  (x => 323, y => 150),
  (x => 324, y => 150),
  (x => 325, y => 150),
  (x => 326, y => 150),
  (x => 327, y => 150),
  (x => 328, y => 150),
  (x => 329, y => 150),
  (x => 330, y => 150),
  (x => 351, y => 150),
  (x => 352, y => 150),
  (x => 353, y => 150),
  (x => 354, y => 150),
  (x => 355, y => 150),
  (x => 356, y => 150),
  (x => 357, y => 150),
  (x => 358, y => 150),
  (x => 365, y => 150),
  (x => 366, y => 150),
  (x => 367, y => 150),
  (x => 368, y => 150),
  (x => 369, y => 150),
  (x => 370, y => 150),
  (x => 381, y => 150),
  (x => 382, y => 150),
  (x => 383, y => 150),
  (x => 384, y => 150),
  (x => 385, y => 150),
  (x => 386, y => 150),
  (x => 387, y => 150),
  (x => 395, y => 150),
  (x => 396, y => 150),
  (x => 397, y => 150),
  (x => 398, y => 150),
  (x => 399, y => 150),
  (x => 400, y => 150),
  (x => 401, y => 150),
  (x => 410, y => 150),
  (x => 411, y => 150),
  (x => 412, y => 150),
  (x => 413, y => 150),
  (x => 414, y => 150),
  (x => 415, y => 150),
  (x => 416, y => 150),
  (x => 424, y => 150),
  (x => 425, y => 150),
  (x => 426, y => 150),
  (x => 427, y => 150),
  (x => 428, y => 150),
  (x => 429, y => 150),
  (x => 430, y => 150),
  (x => 431, y => 150),
  (x => 432, y => 150),
  (x => 433, y => 150),
  (x => 434, y => 150),
  (x => 435, y => 150),
  (x => 439, y => 150),
  (x => 162, y => 151),
  (x => 163, y => 151),
  (x => 164, y => 151),
  (x => 165, y => 151),
  (x => 166, y => 151),
  (x => 167, y => 151),
  (x => 168, y => 151),
  (x => 169, y => 151),
  (x => 179, y => 151),
  (x => 180, y => 151),
  (x => 181, y => 151),
  (x => 182, y => 151),
  (x => 183, y => 151),
  (x => 184, y => 151),
  (x => 185, y => 151),
  (x => 186, y => 151),
  (x => 187, y => 151),
  (x => 188, y => 151),
  (x => 189, y => 151),
  (x => 190, y => 151),
  (x => 191, y => 151),
  (x => 192, y => 151),
  (x => 193, y => 151),
  (x => 216, y => 151),
  (x => 217, y => 151),
  (x => 218, y => 151),
  (x => 219, y => 151),
  (x => 220, y => 151),
  (x => 221, y => 151),
  (x => 222, y => 151),
  (x => 231, y => 151),
  (x => 232, y => 151),
  (x => 233, y => 151),
  (x => 234, y => 151),
  (x => 235, y => 151),
  (x => 236, y => 151),
  (x => 237, y => 151),
  (x => 238, y => 151),
  (x => 239, y => 151),
  (x => 247, y => 151),
  (x => 248, y => 151),
  (x => 249, y => 151),
  (x => 250, y => 151),
  (x => 251, y => 151),
  (x => 252, y => 151),
  (x => 253, y => 151),
  (x => 254, y => 151),
  (x => 255, y => 151),
  (x => 256, y => 151),
  (x => 264, y => 151),
  (x => 265, y => 151),
  (x => 266, y => 151),
  (x => 267, y => 151),
  (x => 268, y => 151),
  (x => 269, y => 151),
  (x => 270, y => 151),
  (x => 271, y => 151),
  (x => 280, y => 151),
  (x => 281, y => 151),
  (x => 282, y => 151),
  (x => 283, y => 151),
  (x => 284, y => 151),
  (x => 285, y => 151),
  (x => 286, y => 151),
  (x => 296, y => 151),
  (x => 297, y => 151),
  (x => 298, y => 151),
  (x => 299, y => 151),
  (x => 300, y => 151),
  (x => 301, y => 151),
  (x => 323, y => 151),
  (x => 324, y => 151),
  (x => 325, y => 151),
  (x => 326, y => 151),
  (x => 327, y => 151),
  (x => 328, y => 151),
  (x => 329, y => 151),
  (x => 330, y => 151),
  (x => 351, y => 151),
  (x => 352, y => 151),
  (x => 353, y => 151),
  (x => 354, y => 151),
  (x => 355, y => 151),
  (x => 356, y => 151),
  (x => 357, y => 151),
  (x => 358, y => 151),
  (x => 365, y => 151),
  (x => 366, y => 151),
  (x => 367, y => 151),
  (x => 368, y => 151),
  (x => 369, y => 151),
  (x => 370, y => 151),
  (x => 371, y => 151),
  (x => 381, y => 151),
  (x => 382, y => 151),
  (x => 383, y => 151),
  (x => 384, y => 151),
  (x => 385, y => 151),
  (x => 386, y => 151),
  (x => 395, y => 151),
  (x => 396, y => 151),
  (x => 397, y => 151),
  (x => 398, y => 151),
  (x => 399, y => 151),
  (x => 400, y => 151),
  (x => 401, y => 151),
  (x => 411, y => 151),
  (x => 412, y => 151),
  (x => 413, y => 151),
  (x => 414, y => 151),
  (x => 415, y => 151),
  (x => 416, y => 151),
  (x => 424, y => 151),
  (x => 425, y => 151),
  (x => 426, y => 151),
  (x => 427, y => 151),
  (x => 428, y => 151),
  (x => 429, y => 151),
  (x => 430, y => 151),
  (x => 431, y => 151),
  (x => 432, y => 151),
  (x => 433, y => 151),
  (x => 162, y => 152),
  (x => 163, y => 152),
  (x => 164, y => 152),
  (x => 165, y => 152),
  (x => 166, y => 152),
  (x => 167, y => 152),
  (x => 168, y => 152),
  (x => 169, y => 152),
  (x => 179, y => 152),
  (x => 180, y => 152),
  (x => 181, y => 152),
  (x => 182, y => 152),
  (x => 183, y => 152),
  (x => 184, y => 152),
  (x => 185, y => 152),
  (x => 186, y => 152),
  (x => 187, y => 152),
  (x => 188, y => 152),
  (x => 189, y => 152),
  (x => 190, y => 152),
  (x => 191, y => 152),
  (x => 192, y => 152),
  (x => 193, y => 152),
  (x => 216, y => 152),
  (x => 217, y => 152),
  (x => 218, y => 152),
  (x => 219, y => 152),
  (x => 220, y => 152),
  (x => 221, y => 152),
  (x => 222, y => 152),
  (x => 231, y => 152),
  (x => 232, y => 152),
  (x => 233, y => 152),
  (x => 234, y => 152),
  (x => 235, y => 152),
  (x => 236, y => 152),
  (x => 237, y => 152),
  (x => 238, y => 152),
  (x => 248, y => 152),
  (x => 249, y => 152),
  (x => 250, y => 152),
  (x => 251, y => 152),
  (x => 252, y => 152),
  (x => 253, y => 152),
  (x => 254, y => 152),
  (x => 255, y => 152),
  (x => 265, y => 152),
  (x => 266, y => 152),
  (x => 267, y => 152),
  (x => 268, y => 152),
  (x => 269, y => 152),
  (x => 270, y => 152),
  (x => 271, y => 152),
  (x => 280, y => 152),
  (x => 281, y => 152),
  (x => 282, y => 152),
  (x => 283, y => 152),
  (x => 284, y => 152),
  (x => 285, y => 152),
  (x => 286, y => 152),
  (x => 297, y => 152),
  (x => 298, y => 152),
  (x => 299, y => 152),
  (x => 300, y => 152),
  (x => 301, y => 152),
  (x => 302, y => 152),
  (x => 323, y => 152),
  (x => 324, y => 152),
  (x => 325, y => 152),
  (x => 326, y => 152),
  (x => 327, y => 152),
  (x => 328, y => 152),
  (x => 329, y => 152),
  (x => 330, y => 152),
  (x => 351, y => 152),
  (x => 352, y => 152),
  (x => 353, y => 152),
  (x => 354, y => 152),
  (x => 355, y => 152),
  (x => 356, y => 152),
  (x => 357, y => 152),
  (x => 358, y => 152),
  (x => 365, y => 152),
  (x => 366, y => 152),
  (x => 367, y => 152),
  (x => 368, y => 152),
  (x => 369, y => 152),
  (x => 370, y => 152),
  (x => 371, y => 152),
  (x => 381, y => 152),
  (x => 382, y => 152),
  (x => 383, y => 152),
  (x => 384, y => 152),
  (x => 385, y => 152),
  (x => 386, y => 152),
  (x => 395, y => 152),
  (x => 396, y => 152),
  (x => 397, y => 152),
  (x => 398, y => 152),
  (x => 399, y => 152),
  (x => 400, y => 152),
  (x => 411, y => 152),
  (x => 412, y => 152),
  (x => 413, y => 152),
  (x => 414, y => 152),
  (x => 415, y => 152),
  (x => 416, y => 152),
  (x => 424, y => 152),
  (x => 425, y => 152),
  (x => 426, y => 152),
  (x => 427, y => 152),
  (x => 428, y => 152),
  (x => 429, y => 152),
  (x => 430, y => 152),
  (x => 431, y => 152),
  (x => 432, y => 152),
  (x => 162, y => 153),
  (x => 163, y => 153),
  (x => 164, y => 153),
  (x => 165, y => 153),
  (x => 166, y => 153),
  (x => 167, y => 153),
  (x => 168, y => 153),
  (x => 169, y => 153),
  (x => 179, y => 153),
  (x => 180, y => 153),
  (x => 181, y => 153),
  (x => 182, y => 153),
  (x => 183, y => 153),
  (x => 184, y => 153),
  (x => 185, y => 153),
  (x => 186, y => 153),
  (x => 187, y => 153),
  (x => 188, y => 153),
  (x => 189, y => 153),
  (x => 190, y => 153),
  (x => 191, y => 153),
  (x => 192, y => 153),
  (x => 193, y => 153),
  (x => 217, y => 153),
  (x => 218, y => 153),
  (x => 219, y => 153),
  (x => 220, y => 153),
  (x => 221, y => 153),
  (x => 222, y => 153),
  (x => 231, y => 153),
  (x => 232, y => 153),
  (x => 233, y => 153),
  (x => 234, y => 153),
  (x => 235, y => 153),
  (x => 236, y => 153),
  (x => 237, y => 153),
  (x => 238, y => 153),
  (x => 248, y => 153),
  (x => 249, y => 153),
  (x => 250, y => 153),
  (x => 251, y => 153),
  (x => 252, y => 153),
  (x => 253, y => 153),
  (x => 254, y => 153),
  (x => 255, y => 153),
  (x => 265, y => 153),
  (x => 266, y => 153),
  (x => 267, y => 153),
  (x => 268, y => 153),
  (x => 269, y => 153),
  (x => 270, y => 153),
  (x => 271, y => 153),
  (x => 280, y => 153),
  (x => 281, y => 153),
  (x => 282, y => 153),
  (x => 283, y => 153),
  (x => 284, y => 153),
  (x => 285, y => 153),
  (x => 297, y => 153),
  (x => 298, y => 153),
  (x => 299, y => 153),
  (x => 300, y => 153),
  (x => 301, y => 153),
  (x => 302, y => 153),
  (x => 323, y => 153),
  (x => 324, y => 153),
  (x => 325, y => 153),
  (x => 326, y => 153),
  (x => 327, y => 153),
  (x => 328, y => 153),
  (x => 329, y => 153),
  (x => 330, y => 153),
  (x => 351, y => 153),
  (x => 352, y => 153),
  (x => 353, y => 153),
  (x => 354, y => 153),
  (x => 355, y => 153),
  (x => 356, y => 153),
  (x => 357, y => 153),
  (x => 358, y => 153),
  (x => 365, y => 153),
  (x => 366, y => 153),
  (x => 367, y => 153),
  (x => 368, y => 153),
  (x => 369, y => 153),
  (x => 370, y => 153),
  (x => 371, y => 153),
  (x => 380, y => 153),
  (x => 381, y => 153),
  (x => 382, y => 153),
  (x => 383, y => 153),
  (x => 384, y => 153),
  (x => 385, y => 153),
  (x => 386, y => 153),
  (x => 394, y => 153),
  (x => 395, y => 153),
  (x => 396, y => 153),
  (x => 397, y => 153),
  (x => 398, y => 153),
  (x => 399, y => 153),
  (x => 400, y => 153),
  (x => 411, y => 153),
  (x => 412, y => 153),
  (x => 413, y => 153),
  (x => 414, y => 153),
  (x => 415, y => 153),
  (x => 416, y => 153),
  (x => 424, y => 153),
  (x => 425, y => 153),
  (x => 426, y => 153),
  (x => 427, y => 153),
  (x => 428, y => 153),
  (x => 429, y => 153),
  (x => 430, y => 153),
  (x => 431, y => 153),
  (x => 432, y => 153),
  (x => 162, y => 154),
  (x => 163, y => 154),
  (x => 164, y => 154),
  (x => 165, y => 154),
  (x => 166, y => 154),
  (x => 167, y => 154),
  (x => 168, y => 154),
  (x => 169, y => 154),
  (x => 179, y => 154),
  (x => 180, y => 154),
  (x => 181, y => 154),
  (x => 182, y => 154),
  (x => 183, y => 154),
  (x => 184, y => 154),
  (x => 185, y => 154),
  (x => 186, y => 154),
  (x => 187, y => 154),
  (x => 188, y => 154),
  (x => 189, y => 154),
  (x => 190, y => 154),
  (x => 191, y => 154),
  (x => 192, y => 154),
  (x => 193, y => 154),
  (x => 217, y => 154),
  (x => 218, y => 154),
  (x => 219, y => 154),
  (x => 220, y => 154),
  (x => 221, y => 154),
  (x => 222, y => 154),
  (x => 231, y => 154),
  (x => 232, y => 154),
  (x => 233, y => 154),
  (x => 234, y => 154),
  (x => 235, y => 154),
  (x => 236, y => 154),
  (x => 237, y => 154),
  (x => 248, y => 154),
  (x => 249, y => 154),
  (x => 250, y => 154),
  (x => 251, y => 154),
  (x => 252, y => 154),
  (x => 253, y => 154),
  (x => 254, y => 154),
  (x => 255, y => 154),
  (x => 265, y => 154),
  (x => 266, y => 154),
  (x => 267, y => 154),
  (x => 268, y => 154),
  (x => 269, y => 154),
  (x => 270, y => 154),
  (x => 271, y => 154),
  (x => 280, y => 154),
  (x => 281, y => 154),
  (x => 282, y => 154),
  (x => 283, y => 154),
  (x => 284, y => 154),
  (x => 285, y => 154),
  (x => 297, y => 154),
  (x => 298, y => 154),
  (x => 299, y => 154),
  (x => 300, y => 154),
  (x => 301, y => 154),
  (x => 302, y => 154),
  (x => 323, y => 154),
  (x => 324, y => 154),
  (x => 325, y => 154),
  (x => 326, y => 154),
  (x => 327, y => 154),
  (x => 328, y => 154),
  (x => 329, y => 154),
  (x => 330, y => 154),
  (x => 351, y => 154),
  (x => 352, y => 154),
  (x => 353, y => 154),
  (x => 354, y => 154),
  (x => 355, y => 154),
  (x => 356, y => 154),
  (x => 357, y => 154),
  (x => 358, y => 154),
  (x => 366, y => 154),
  (x => 367, y => 154),
  (x => 368, y => 154),
  (x => 369, y => 154),
  (x => 370, y => 154),
  (x => 371, y => 154),
  (x => 380, y => 154),
  (x => 381, y => 154),
  (x => 382, y => 154),
  (x => 383, y => 154),
  (x => 384, y => 154),
  (x => 385, y => 154),
  (x => 386, y => 154),
  (x => 394, y => 154),
  (x => 395, y => 154),
  (x => 396, y => 154),
  (x => 397, y => 154),
  (x => 398, y => 154),
  (x => 399, y => 154),
  (x => 400, y => 154),
  (x => 411, y => 154),
  (x => 412, y => 154),
  (x => 413, y => 154),
  (x => 414, y => 154),
  (x => 415, y => 154),
  (x => 416, y => 154),
  (x => 417, y => 154),
  (x => 424, y => 154),
  (x => 425, y => 154),
  (x => 426, y => 154),
  (x => 427, y => 154),
  (x => 428, y => 154),
  (x => 429, y => 154),
  (x => 430, y => 154),
  (x => 431, y => 154),
  (x => 162, y => 155),
  (x => 163, y => 155),
  (x => 164, y => 155),
  (x => 165, y => 155),
  (x => 166, y => 155),
  (x => 167, y => 155),
  (x => 168, y => 155),
  (x => 169, y => 155),
  (x => 179, y => 155),
  (x => 180, y => 155),
  (x => 181, y => 155),
  (x => 182, y => 155),
  (x => 183, y => 155),
  (x => 184, y => 155),
  (x => 185, y => 155),
  (x => 186, y => 155),
  (x => 187, y => 155),
  (x => 188, y => 155),
  (x => 189, y => 155),
  (x => 190, y => 155),
  (x => 191, y => 155),
  (x => 192, y => 155),
  (x => 193, y => 155),
  (x => 216, y => 155),
  (x => 217, y => 155),
  (x => 218, y => 155),
  (x => 219, y => 155),
  (x => 220, y => 155),
  (x => 221, y => 155),
  (x => 222, y => 155),
  (x => 231, y => 155),
  (x => 232, y => 155),
  (x => 233, y => 155),
  (x => 234, y => 155),
  (x => 235, y => 155),
  (x => 236, y => 155),
  (x => 237, y => 155),
  (x => 248, y => 155),
  (x => 249, y => 155),
  (x => 250, y => 155),
  (x => 251, y => 155),
  (x => 252, y => 155),
  (x => 253, y => 155),
  (x => 254, y => 155),
  (x => 266, y => 155),
  (x => 267, y => 155),
  (x => 268, y => 155),
  (x => 269, y => 155),
  (x => 270, y => 155),
  (x => 271, y => 155),
  (x => 272, y => 155),
  (x => 279, y => 155),
  (x => 280, y => 155),
  (x => 281, y => 155),
  (x => 282, y => 155),
  (x => 283, y => 155),
  (x => 284, y => 155),
  (x => 285, y => 155),
  (x => 297, y => 155),
  (x => 298, y => 155),
  (x => 299, y => 155),
  (x => 300, y => 155),
  (x => 301, y => 155),
  (x => 302, y => 155),
  (x => 323, y => 155),
  (x => 324, y => 155),
  (x => 325, y => 155),
  (x => 326, y => 155),
  (x => 327, y => 155),
  (x => 328, y => 155),
  (x => 329, y => 155),
  (x => 330, y => 155),
  (x => 351, y => 155),
  (x => 352, y => 155),
  (x => 353, y => 155),
  (x => 354, y => 155),
  (x => 355, y => 155),
  (x => 356, y => 155),
  (x => 357, y => 155),
  (x => 358, y => 155),
  (x => 366, y => 155),
  (x => 367, y => 155),
  (x => 368, y => 155),
  (x => 369, y => 155),
  (x => 370, y => 155),
  (x => 371, y => 155),
  (x => 372, y => 155),
  (x => 380, y => 155),
  (x => 381, y => 155),
  (x => 382, y => 155),
  (x => 383, y => 155),
  (x => 384, y => 155),
  (x => 385, y => 155),
  (x => 394, y => 155),
  (x => 395, y => 155),
  (x => 396, y => 155),
  (x => 397, y => 155),
  (x => 398, y => 155),
  (x => 399, y => 155),
  (x => 412, y => 155),
  (x => 413, y => 155),
  (x => 414, y => 155),
  (x => 415, y => 155),
  (x => 416, y => 155),
  (x => 417, y => 155),
  (x => 424, y => 155),
  (x => 425, y => 155),
  (x => 426, y => 155),
  (x => 427, y => 155),
  (x => 428, y => 155),
  (x => 429, y => 155),
  (x => 430, y => 155),
  (x => 431, y => 155),
  (x => 162, y => 156),
  (x => 163, y => 156),
  (x => 164, y => 156),
  (x => 165, y => 156),
  (x => 166, y => 156),
  (x => 167, y => 156),
  (x => 168, y => 156),
  (x => 169, y => 156),
  (x => 179, y => 156),
  (x => 180, y => 156),
  (x => 181, y => 156),
  (x => 182, y => 156),
  (x => 183, y => 156),
  (x => 184, y => 156),
  (x => 185, y => 156),
  (x => 186, y => 156),
  (x => 187, y => 156),
  (x => 188, y => 156),
  (x => 189, y => 156),
  (x => 190, y => 156),
  (x => 191, y => 156),
  (x => 192, y => 156),
  (x => 193, y => 156),
  (x => 212, y => 156),
  (x => 213, y => 156),
  (x => 214, y => 156),
  (x => 215, y => 156),
  (x => 216, y => 156),
  (x => 217, y => 156),
  (x => 218, y => 156),
  (x => 219, y => 156),
  (x => 220, y => 156),
  (x => 221, y => 156),
  (x => 222, y => 156),
  (x => 231, y => 156),
  (x => 232, y => 156),
  (x => 233, y => 156),
  (x => 234, y => 156),
  (x => 235, y => 156),
  (x => 236, y => 156),
  (x => 237, y => 156),
  (x => 248, y => 156),
  (x => 249, y => 156),
  (x => 250, y => 156),
  (x => 251, y => 156),
  (x => 252, y => 156),
  (x => 253, y => 156),
  (x => 254, y => 156),
  (x => 266, y => 156),
  (x => 267, y => 156),
  (x => 268, y => 156),
  (x => 269, y => 156),
  (x => 270, y => 156),
  (x => 271, y => 156),
  (x => 272, y => 156),
  (x => 279, y => 156),
  (x => 280, y => 156),
  (x => 281, y => 156),
  (x => 282, y => 156),
  (x => 283, y => 156),
  (x => 284, y => 156),
  (x => 285, y => 156),
  (x => 297, y => 156),
  (x => 298, y => 156),
  (x => 299, y => 156),
  (x => 300, y => 156),
  (x => 301, y => 156),
  (x => 302, y => 156),
  (x => 323, y => 156),
  (x => 324, y => 156),
  (x => 325, y => 156),
  (x => 326, y => 156),
  (x => 327, y => 156),
  (x => 328, y => 156),
  (x => 329, y => 156),
  (x => 330, y => 156),
  (x => 351, y => 156),
  (x => 352, y => 156),
  (x => 353, y => 156),
  (x => 354, y => 156),
  (x => 355, y => 156),
  (x => 356, y => 156),
  (x => 357, y => 156),
  (x => 358, y => 156),
  (x => 366, y => 156),
  (x => 367, y => 156),
  (x => 368, y => 156),
  (x => 369, y => 156),
  (x => 370, y => 156),
  (x => 371, y => 156),
  (x => 372, y => 156),
  (x => 380, y => 156),
  (x => 381, y => 156),
  (x => 382, y => 156),
  (x => 383, y => 156),
  (x => 384, y => 156),
  (x => 385, y => 156),
  (x => 394, y => 156),
  (x => 395, y => 156),
  (x => 396, y => 156),
  (x => 397, y => 156),
  (x => 398, y => 156),
  (x => 399, y => 156),
  (x => 412, y => 156),
  (x => 413, y => 156),
  (x => 414, y => 156),
  (x => 415, y => 156),
  (x => 416, y => 156),
  (x => 417, y => 156),
  (x => 424, y => 156),
  (x => 425, y => 156),
  (x => 426, y => 156),
  (x => 427, y => 156),
  (x => 428, y => 156),
  (x => 429, y => 156),
  (x => 430, y => 156),
  (x => 431, y => 156),
  (x => 162, y => 157),
  (x => 163, y => 157),
  (x => 164, y => 157),
  (x => 165, y => 157),
  (x => 166, y => 157),
  (x => 167, y => 157),
  (x => 168, y => 157),
  (x => 169, y => 157),
  (x => 179, y => 157),
  (x => 180, y => 157),
  (x => 181, y => 157),
  (x => 182, y => 157),
  (x => 183, y => 157),
  (x => 184, y => 157),
  (x => 185, y => 157),
  (x => 186, y => 157),
  (x => 187, y => 157),
  (x => 188, y => 157),
  (x => 189, y => 157),
  (x => 190, y => 157),
  (x => 191, y => 157),
  (x => 192, y => 157),
  (x => 193, y => 157),
  (x => 207, y => 157),
  (x => 208, y => 157),
  (x => 209, y => 157),
  (x => 210, y => 157),
  (x => 211, y => 157),
  (x => 212, y => 157),
  (x => 213, y => 157),
  (x => 214, y => 157),
  (x => 215, y => 157),
  (x => 216, y => 157),
  (x => 217, y => 157),
  (x => 218, y => 157),
  (x => 219, y => 157),
  (x => 220, y => 157),
  (x => 221, y => 157),
  (x => 222, y => 157),
  (x => 231, y => 157),
  (x => 232, y => 157),
  (x => 233, y => 157),
  (x => 234, y => 157),
  (x => 235, y => 157),
  (x => 236, y => 157),
  (x => 237, y => 157),
  (x => 248, y => 157),
  (x => 249, y => 157),
  (x => 250, y => 157),
  (x => 251, y => 157),
  (x => 252, y => 157),
  (x => 253, y => 157),
  (x => 254, y => 157),
  (x => 266, y => 157),
  (x => 267, y => 157),
  (x => 268, y => 157),
  (x => 269, y => 157),
  (x => 270, y => 157),
  (x => 271, y => 157),
  (x => 272, y => 157),
  (x => 279, y => 157),
  (x => 280, y => 157),
  (x => 281, y => 157),
  (x => 282, y => 157),
  (x => 283, y => 157),
  (x => 284, y => 157),
  (x => 285, y => 157),
  (x => 297, y => 157),
  (x => 298, y => 157),
  (x => 299, y => 157),
  (x => 300, y => 157),
  (x => 301, y => 157),
  (x => 302, y => 157),
  (x => 323, y => 157),
  (x => 324, y => 157),
  (x => 325, y => 157),
  (x => 326, y => 157),
  (x => 327, y => 157),
  (x => 328, y => 157),
  (x => 329, y => 157),
  (x => 330, y => 157),
  (x => 351, y => 157),
  (x => 352, y => 157),
  (x => 353, y => 157),
  (x => 354, y => 157),
  (x => 355, y => 157),
  (x => 356, y => 157),
  (x => 357, y => 157),
  (x => 358, y => 157),
  (x => 366, y => 157),
  (x => 367, y => 157),
  (x => 368, y => 157),
  (x => 369, y => 157),
  (x => 370, y => 157),
  (x => 371, y => 157),
  (x => 372, y => 157),
  (x => 380, y => 157),
  (x => 381, y => 157),
  (x => 382, y => 157),
  (x => 383, y => 157),
  (x => 384, y => 157),
  (x => 385, y => 157),
  (x => 394, y => 157),
  (x => 395, y => 157),
  (x => 396, y => 157),
  (x => 397, y => 157),
  (x => 398, y => 157),
  (x => 399, y => 157),
  (x => 412, y => 157),
  (x => 413, y => 157),
  (x => 414, y => 157),
  (x => 415, y => 157),
  (x => 416, y => 157),
  (x => 417, y => 157),
  (x => 424, y => 157),
  (x => 425, y => 157),
  (x => 426, y => 157),
  (x => 427, y => 157),
  (x => 428, y => 157),
  (x => 429, y => 157),
  (x => 430, y => 157),
  (x => 162, y => 158),
  (x => 163, y => 158),
  (x => 164, y => 158),
  (x => 165, y => 158),
  (x => 166, y => 158),
  (x => 167, y => 158),
  (x => 168, y => 158),
  (x => 169, y => 158),
  (x => 187, y => 158),
  (x => 188, y => 158),
  (x => 189, y => 158),
  (x => 190, y => 158),
  (x => 191, y => 158),
  (x => 192, y => 158),
  (x => 193, y => 158),
  (x => 205, y => 158),
  (x => 206, y => 158),
  (x => 207, y => 158),
  (x => 208, y => 158),
  (x => 209, y => 158),
  (x => 210, y => 158),
  (x => 211, y => 158),
  (x => 212, y => 158),
  (x => 213, y => 158),
  (x => 214, y => 158),
  (x => 215, y => 158),
  (x => 216, y => 158),
  (x => 217, y => 158),
  (x => 218, y => 158),
  (x => 219, y => 158),
  (x => 220, y => 158),
  (x => 221, y => 158),
  (x => 222, y => 158),
  (x => 231, y => 158),
  (x => 232, y => 158),
  (x => 233, y => 158),
  (x => 234, y => 158),
  (x => 235, y => 158),
  (x => 236, y => 158),
  (x => 237, y => 158),
  (x => 248, y => 158),
  (x => 249, y => 158),
  (x => 250, y => 158),
  (x => 251, y => 158),
  (x => 252, y => 158),
  (x => 253, y => 158),
  (x => 254, y => 158),
  (x => 266, y => 158),
  (x => 267, y => 158),
  (x => 268, y => 158),
  (x => 269, y => 158),
  (x => 270, y => 158),
  (x => 271, y => 158),
  (x => 272, y => 158),
  (x => 279, y => 158),
  (x => 280, y => 158),
  (x => 281, y => 158),
  (x => 282, y => 158),
  (x => 283, y => 158),
  (x => 284, y => 158),
  (x => 285, y => 158),
  (x => 286, y => 158),
  (x => 287, y => 158),
  (x => 288, y => 158),
  (x => 289, y => 158),
  (x => 290, y => 158),
  (x => 291, y => 158),
  (x => 292, y => 158),
  (x => 293, y => 158),
  (x => 294, y => 158),
  (x => 295, y => 158),
  (x => 296, y => 158),
  (x => 297, y => 158),
  (x => 298, y => 158),
  (x => 299, y => 158),
  (x => 300, y => 158),
  (x => 301, y => 158),
  (x => 302, y => 158),
  (x => 323, y => 158),
  (x => 324, y => 158),
  (x => 325, y => 158),
  (x => 326, y => 158),
  (x => 327, y => 158),
  (x => 328, y => 158),
  (x => 329, y => 158),
  (x => 330, y => 158),
  (x => 351, y => 158),
  (x => 352, y => 158),
  (x => 353, y => 158),
  (x => 354, y => 158),
  (x => 355, y => 158),
  (x => 356, y => 158),
  (x => 357, y => 158),
  (x => 358, y => 158),
  (x => 367, y => 158),
  (x => 368, y => 158),
  (x => 369, y => 158),
  (x => 370, y => 158),
  (x => 371, y => 158),
  (x => 372, y => 158),
  (x => 379, y => 158),
  (x => 380, y => 158),
  (x => 381, y => 158),
  (x => 382, y => 158),
  (x => 383, y => 158),
  (x => 384, y => 158),
  (x => 385, y => 158),
  (x => 394, y => 158),
  (x => 395, y => 158),
  (x => 396, y => 158),
  (x => 397, y => 158),
  (x => 398, y => 158),
  (x => 399, y => 158),
  (x => 400, y => 158),
  (x => 401, y => 158),
  (x => 402, y => 158),
  (x => 403, y => 158),
  (x => 404, y => 158),
  (x => 405, y => 158),
  (x => 406, y => 158),
  (x => 407, y => 158),
  (x => 408, y => 158),
  (x => 409, y => 158),
  (x => 410, y => 158),
  (x => 411, y => 158),
  (x => 412, y => 158),
  (x => 413, y => 158),
  (x => 414, y => 158),
  (x => 415, y => 158),
  (x => 416, y => 158),
  (x => 417, y => 158),
  (x => 424, y => 158),
  (x => 425, y => 158),
  (x => 426, y => 158),
  (x => 427, y => 158),
  (x => 428, y => 158),
  (x => 429, y => 158),
  (x => 430, y => 158),
  (x => 162, y => 159),
  (x => 163, y => 159),
  (x => 164, y => 159),
  (x => 165, y => 159),
  (x => 166, y => 159),
  (x => 167, y => 159),
  (x => 168, y => 159),
  (x => 169, y => 159),
  (x => 187, y => 159),
  (x => 188, y => 159),
  (x => 189, y => 159),
  (x => 190, y => 159),
  (x => 191, y => 159),
  (x => 192, y => 159),
  (x => 193, y => 159),
  (x => 203, y => 159),
  (x => 204, y => 159),
  (x => 205, y => 159),
  (x => 206, y => 159),
  (x => 207, y => 159),
  (x => 208, y => 159),
  (x => 209, y => 159),
  (x => 210, y => 159),
  (x => 211, y => 159),
  (x => 212, y => 159),
  (x => 213, y => 159),
  (x => 214, y => 159),
  (x => 215, y => 159),
  (x => 216, y => 159),
  (x => 217, y => 159),
  (x => 218, y => 159),
  (x => 219, y => 159),
  (x => 220, y => 159),
  (x => 221, y => 159),
  (x => 222, y => 159),
  (x => 231, y => 159),
  (x => 232, y => 159),
  (x => 233, y => 159),
  (x => 234, y => 159),
  (x => 235, y => 159),
  (x => 236, y => 159),
  (x => 237, y => 159),
  (x => 248, y => 159),
  (x => 249, y => 159),
  (x => 250, y => 159),
  (x => 251, y => 159),
  (x => 252, y => 159),
  (x => 253, y => 159),
  (x => 254, y => 159),
  (x => 266, y => 159),
  (x => 267, y => 159),
  (x => 268, y => 159),
  (x => 269, y => 159),
  (x => 270, y => 159),
  (x => 271, y => 159),
  (x => 272, y => 159),
  (x => 279, y => 159),
  (x => 280, y => 159),
  (x => 281, y => 159),
  (x => 282, y => 159),
  (x => 283, y => 159),
  (x => 284, y => 159),
  (x => 285, y => 159),
  (x => 286, y => 159),
  (x => 287, y => 159),
  (x => 288, y => 159),
  (x => 289, y => 159),
  (x => 290, y => 159),
  (x => 291, y => 159),
  (x => 292, y => 159),
  (x => 293, y => 159),
  (x => 294, y => 159),
  (x => 295, y => 159),
  (x => 296, y => 159),
  (x => 297, y => 159),
  (x => 298, y => 159),
  (x => 299, y => 159),
  (x => 300, y => 159),
  (x => 301, y => 159),
  (x => 302, y => 159),
  (x => 324, y => 159),
  (x => 325, y => 159),
  (x => 326, y => 159),
  (x => 327, y => 159),
  (x => 328, y => 159),
  (x => 329, y => 159),
  (x => 330, y => 159),
  (x => 351, y => 159),
  (x => 352, y => 159),
  (x => 353, y => 159),
  (x => 354, y => 159),
  (x => 355, y => 159),
  (x => 356, y => 159),
  (x => 357, y => 159),
  (x => 367, y => 159),
  (x => 368, y => 159),
  (x => 369, y => 159),
  (x => 370, y => 159),
  (x => 371, y => 159),
  (x => 372, y => 159),
  (x => 379, y => 159),
  (x => 380, y => 159),
  (x => 381, y => 159),
  (x => 382, y => 159),
  (x => 383, y => 159),
  (x => 384, y => 159),
  (x => 393, y => 159),
  (x => 394, y => 159),
  (x => 395, y => 159),
  (x => 396, y => 159),
  (x => 397, y => 159),
  (x => 398, y => 159),
  (x => 399, y => 159),
  (x => 400, y => 159),
  (x => 401, y => 159),
  (x => 402, y => 159),
  (x => 403, y => 159),
  (x => 404, y => 159),
  (x => 405, y => 159),
  (x => 406, y => 159),
  (x => 407, y => 159),
  (x => 408, y => 159),
  (x => 409, y => 159),
  (x => 410, y => 159),
  (x => 411, y => 159),
  (x => 412, y => 159),
  (x => 413, y => 159),
  (x => 414, y => 159),
  (x => 415, y => 159),
  (x => 416, y => 159),
  (x => 417, y => 159),
  (x => 424, y => 159),
  (x => 425, y => 159),
  (x => 426, y => 159),
  (x => 427, y => 159),
  (x => 428, y => 159),
  (x => 429, y => 159),
  (x => 430, y => 159),
  (x => 163, y => 160),
  (x => 164, y => 160),
  (x => 165, y => 160),
  (x => 166, y => 160),
  (x => 167, y => 160),
  (x => 168, y => 160),
  (x => 169, y => 160),
  (x => 187, y => 160),
  (x => 188, y => 160),
  (x => 189, y => 160),
  (x => 190, y => 160),
  (x => 191, y => 160),
  (x => 192, y => 160),
  (x => 193, y => 160),
  (x => 202, y => 160),
  (x => 203, y => 160),
  (x => 204, y => 160),
  (x => 205, y => 160),
  (x => 206, y => 160),
  (x => 207, y => 160),
  (x => 208, y => 160),
  (x => 209, y => 160),
  (x => 210, y => 160),
  (x => 211, y => 160),
  (x => 212, y => 160),
  (x => 213, y => 160),
  (x => 214, y => 160),
  (x => 215, y => 160),
  (x => 216, y => 160),
  (x => 217, y => 160),
  (x => 218, y => 160),
  (x => 219, y => 160),
  (x => 220, y => 160),
  (x => 221, y => 160),
  (x => 222, y => 160),
  (x => 231, y => 160),
  (x => 232, y => 160),
  (x => 233, y => 160),
  (x => 234, y => 160),
  (x => 235, y => 160),
  (x => 236, y => 160),
  (x => 237, y => 160),
  (x => 248, y => 160),
  (x => 249, y => 160),
  (x => 250, y => 160),
  (x => 251, y => 160),
  (x => 252, y => 160),
  (x => 253, y => 160),
  (x => 254, y => 160),
  (x => 266, y => 160),
  (x => 267, y => 160),
  (x => 268, y => 160),
  (x => 269, y => 160),
  (x => 270, y => 160),
  (x => 271, y => 160),
  (x => 272, y => 160),
  (x => 279, y => 160),
  (x => 280, y => 160),
  (x => 281, y => 160),
  (x => 282, y => 160),
  (x => 283, y => 160),
  (x => 284, y => 160),
  (x => 285, y => 160),
  (x => 286, y => 160),
  (x => 287, y => 160),
  (x => 288, y => 160),
  (x => 289, y => 160),
  (x => 290, y => 160),
  (x => 291, y => 160),
  (x => 292, y => 160),
  (x => 293, y => 160),
  (x => 294, y => 160),
  (x => 295, y => 160),
  (x => 296, y => 160),
  (x => 297, y => 160),
  (x => 298, y => 160),
  (x => 299, y => 160),
  (x => 300, y => 160),
  (x => 301, y => 160),
  (x => 302, y => 160),
  (x => 324, y => 160),
  (x => 325, y => 160),
  (x => 326, y => 160),
  (x => 327, y => 160),
  (x => 328, y => 160),
  (x => 329, y => 160),
  (x => 330, y => 160),
  (x => 331, y => 160),
  (x => 351, y => 160),
  (x => 352, y => 160),
  (x => 353, y => 160),
  (x => 354, y => 160),
  (x => 355, y => 160),
  (x => 356, y => 160),
  (x => 357, y => 160),
  (x => 367, y => 160),
  (x => 368, y => 160),
  (x => 369, y => 160),
  (x => 370, y => 160),
  (x => 371, y => 160),
  (x => 372, y => 160),
  (x => 373, y => 160),
  (x => 379, y => 160),
  (x => 380, y => 160),
  (x => 381, y => 160),
  (x => 382, y => 160),
  (x => 383, y => 160),
  (x => 384, y => 160),
  (x => 393, y => 160),
  (x => 394, y => 160),
  (x => 395, y => 160),
  (x => 396, y => 160),
  (x => 397, y => 160),
  (x => 398, y => 160),
  (x => 399, y => 160),
  (x => 400, y => 160),
  (x => 401, y => 160),
  (x => 402, y => 160),
  (x => 403, y => 160),
  (x => 404, y => 160),
  (x => 405, y => 160),
  (x => 406, y => 160),
  (x => 407, y => 160),
  (x => 408, y => 160),
  (x => 409, y => 160),
  (x => 410, y => 160),
  (x => 411, y => 160),
  (x => 412, y => 160),
  (x => 413, y => 160),
  (x => 414, y => 160),
  (x => 415, y => 160),
  (x => 416, y => 160),
  (x => 417, y => 160),
  (x => 424, y => 160),
  (x => 425, y => 160),
  (x => 426, y => 160),
  (x => 427, y => 160),
  (x => 428, y => 160),
  (x => 429, y => 160),
  (x => 430, y => 160),
  (x => 163, y => 161),
  (x => 164, y => 161),
  (x => 165, y => 161),
  (x => 166, y => 161),
  (x => 167, y => 161),
  (x => 168, y => 161),
  (x => 169, y => 161),
  (x => 170, y => 161),
  (x => 187, y => 161),
  (x => 188, y => 161),
  (x => 189, y => 161),
  (x => 190, y => 161),
  (x => 191, y => 161),
  (x => 192, y => 161),
  (x => 193, y => 161),
  (x => 202, y => 161),
  (x => 203, y => 161),
  (x => 204, y => 161),
  (x => 205, y => 161),
  (x => 206, y => 161),
  (x => 207, y => 161),
  (x => 208, y => 161),
  (x => 209, y => 161),
  (x => 210, y => 161),
  (x => 217, y => 161),
  (x => 218, y => 161),
  (x => 219, y => 161),
  (x => 220, y => 161),
  (x => 221, y => 161),
  (x => 222, y => 161),
  (x => 231, y => 161),
  (x => 232, y => 161),
  (x => 233, y => 161),
  (x => 234, y => 161),
  (x => 235, y => 161),
  (x => 236, y => 161),
  (x => 237, y => 161),
  (x => 248, y => 161),
  (x => 249, y => 161),
  (x => 250, y => 161),
  (x => 251, y => 161),
  (x => 252, y => 161),
  (x => 253, y => 161),
  (x => 254, y => 161),
  (x => 266, y => 161),
  (x => 267, y => 161),
  (x => 268, y => 161),
  (x => 269, y => 161),
  (x => 270, y => 161),
  (x => 271, y => 161),
  (x => 272, y => 161),
  (x => 279, y => 161),
  (x => 280, y => 161),
  (x => 281, y => 161),
  (x => 282, y => 161),
  (x => 283, y => 161),
  (x => 284, y => 161),
  (x => 285, y => 161),
  (x => 286, y => 161),
  (x => 287, y => 161),
  (x => 288, y => 161),
  (x => 289, y => 161),
  (x => 290, y => 161),
  (x => 291, y => 161),
  (x => 292, y => 161),
  (x => 293, y => 161),
  (x => 294, y => 161),
  (x => 295, y => 161),
  (x => 296, y => 161),
  (x => 297, y => 161),
  (x => 298, y => 161),
  (x => 299, y => 161),
  (x => 300, y => 161),
  (x => 301, y => 161),
  (x => 302, y => 161),
  (x => 324, y => 161),
  (x => 325, y => 161),
  (x => 326, y => 161),
  (x => 327, y => 161),
  (x => 328, y => 161),
  (x => 329, y => 161),
  (x => 330, y => 161),
  (x => 331, y => 161),
  (x => 350, y => 161),
  (x => 351, y => 161),
  (x => 352, y => 161),
  (x => 353, y => 161),
  (x => 354, y => 161),
  (x => 355, y => 161),
  (x => 356, y => 161),
  (x => 357, y => 161),
  (x => 367, y => 161),
  (x => 368, y => 161),
  (x => 369, y => 161),
  (x => 370, y => 161),
  (x => 371, y => 161),
  (x => 372, y => 161),
  (x => 373, y => 161),
  (x => 379, y => 161),
  (x => 380, y => 161),
  (x => 381, y => 161),
  (x => 382, y => 161),
  (x => 383, y => 161),
  (x => 384, y => 161),
  (x => 393, y => 161),
  (x => 394, y => 161),
  (x => 395, y => 161),
  (x => 396, y => 161),
  (x => 397, y => 161),
  (x => 398, y => 161),
  (x => 399, y => 161),
  (x => 400, y => 161),
  (x => 401, y => 161),
  (x => 402, y => 161),
  (x => 403, y => 161),
  (x => 404, y => 161),
  (x => 405, y => 161),
  (x => 406, y => 161),
  (x => 407, y => 161),
  (x => 408, y => 161),
  (x => 409, y => 161),
  (x => 410, y => 161),
  (x => 411, y => 161),
  (x => 412, y => 161),
  (x => 413, y => 161),
  (x => 414, y => 161),
  (x => 415, y => 161),
  (x => 416, y => 161),
  (x => 417, y => 161),
  (x => 424, y => 161),
  (x => 425, y => 161),
  (x => 426, y => 161),
  (x => 427, y => 161),
  (x => 428, y => 161),
  (x => 429, y => 161),
  (x => 430, y => 161),
  (x => 163, y => 162),
  (x => 164, y => 162),
  (x => 165, y => 162),
  (x => 166, y => 162),
  (x => 167, y => 162),
  (x => 168, y => 162),
  (x => 169, y => 162),
  (x => 170, y => 162),
  (x => 187, y => 162),
  (x => 188, y => 162),
  (x => 189, y => 162),
  (x => 190, y => 162),
  (x => 191, y => 162),
  (x => 192, y => 162),
  (x => 193, y => 162),
  (x => 201, y => 162),
  (x => 202, y => 162),
  (x => 203, y => 162),
  (x => 204, y => 162),
  (x => 205, y => 162),
  (x => 206, y => 162),
  (x => 207, y => 162),
  (x => 208, y => 162),
  (x => 217, y => 162),
  (x => 218, y => 162),
  (x => 219, y => 162),
  (x => 220, y => 162),
  (x => 221, y => 162),
  (x => 222, y => 162),
  (x => 231, y => 162),
  (x => 232, y => 162),
  (x => 233, y => 162),
  (x => 234, y => 162),
  (x => 235, y => 162),
  (x => 236, y => 162),
  (x => 237, y => 162),
  (x => 248, y => 162),
  (x => 249, y => 162),
  (x => 250, y => 162),
  (x => 251, y => 162),
  (x => 252, y => 162),
  (x => 253, y => 162),
  (x => 254, y => 162),
  (x => 266, y => 162),
  (x => 267, y => 162),
  (x => 268, y => 162),
  (x => 269, y => 162),
  (x => 270, y => 162),
  (x => 271, y => 162),
  (x => 272, y => 162),
  (x => 279, y => 162),
  (x => 280, y => 162),
  (x => 281, y => 162),
  (x => 282, y => 162),
  (x => 283, y => 162),
  (x => 284, y => 162),
  (x => 285, y => 162),
  (x => 286, y => 162),
  (x => 287, y => 162),
  (x => 288, y => 162),
  (x => 289, y => 162),
  (x => 290, y => 162),
  (x => 291, y => 162),
  (x => 292, y => 162),
  (x => 293, y => 162),
  (x => 294, y => 162),
  (x => 295, y => 162),
  (x => 296, y => 162),
  (x => 297, y => 162),
  (x => 298, y => 162),
  (x => 299, y => 162),
  (x => 300, y => 162),
  (x => 301, y => 162),
  (x => 302, y => 162),
  (x => 324, y => 162),
  (x => 325, y => 162),
  (x => 326, y => 162),
  (x => 327, y => 162),
  (x => 328, y => 162),
  (x => 329, y => 162),
  (x => 330, y => 162),
  (x => 331, y => 162),
  (x => 350, y => 162),
  (x => 351, y => 162),
  (x => 352, y => 162),
  (x => 353, y => 162),
  (x => 354, y => 162),
  (x => 355, y => 162),
  (x => 356, y => 162),
  (x => 357, y => 162),
  (x => 368, y => 162),
  (x => 369, y => 162),
  (x => 370, y => 162),
  (x => 371, y => 162),
  (x => 372, y => 162),
  (x => 373, y => 162),
  (x => 378, y => 162),
  (x => 379, y => 162),
  (x => 380, y => 162),
  (x => 381, y => 162),
  (x => 382, y => 162),
  (x => 383, y => 162),
  (x => 393, y => 162),
  (x => 394, y => 162),
  (x => 395, y => 162),
  (x => 396, y => 162),
  (x => 397, y => 162),
  (x => 398, y => 162),
  (x => 399, y => 162),
  (x => 400, y => 162),
  (x => 401, y => 162),
  (x => 402, y => 162),
  (x => 403, y => 162),
  (x => 404, y => 162),
  (x => 405, y => 162),
  (x => 406, y => 162),
  (x => 407, y => 162),
  (x => 408, y => 162),
  (x => 409, y => 162),
  (x => 410, y => 162),
  (x => 411, y => 162),
  (x => 412, y => 162),
  (x => 413, y => 162),
  (x => 414, y => 162),
  (x => 415, y => 162),
  (x => 416, y => 162),
  (x => 417, y => 162),
  (x => 424, y => 162),
  (x => 425, y => 162),
  (x => 426, y => 162),
  (x => 427, y => 162),
  (x => 428, y => 162),
  (x => 429, y => 162),
  (x => 430, y => 162),
  (x => 163, y => 163),
  (x => 164, y => 163),
  (x => 165, y => 163),
  (x => 166, y => 163),
  (x => 167, y => 163),
  (x => 168, y => 163),
  (x => 169, y => 163),
  (x => 170, y => 163),
  (x => 187, y => 163),
  (x => 188, y => 163),
  (x => 189, y => 163),
  (x => 190, y => 163),
  (x => 191, y => 163),
  (x => 192, y => 163),
  (x => 193, y => 163),
  (x => 201, y => 163),
  (x => 202, y => 163),
  (x => 203, y => 163),
  (x => 204, y => 163),
  (x => 205, y => 163),
  (x => 206, y => 163),
  (x => 217, y => 163),
  (x => 218, y => 163),
  (x => 219, y => 163),
  (x => 220, y => 163),
  (x => 221, y => 163),
  (x => 222, y => 163),
  (x => 231, y => 163),
  (x => 232, y => 163),
  (x => 233, y => 163),
  (x => 234, y => 163),
  (x => 235, y => 163),
  (x => 236, y => 163),
  (x => 237, y => 163),
  (x => 248, y => 163),
  (x => 249, y => 163),
  (x => 250, y => 163),
  (x => 251, y => 163),
  (x => 252, y => 163),
  (x => 253, y => 163),
  (x => 254, y => 163),
  (x => 266, y => 163),
  (x => 267, y => 163),
  (x => 268, y => 163),
  (x => 269, y => 163),
  (x => 270, y => 163),
  (x => 271, y => 163),
  (x => 272, y => 163),
  (x => 279, y => 163),
  (x => 280, y => 163),
  (x => 281, y => 163),
  (x => 282, y => 163),
  (x => 283, y => 163),
  (x => 284, y => 163),
  (x => 285, y => 163),
  (x => 324, y => 163),
  (x => 325, y => 163),
  (x => 326, y => 163),
  (x => 327, y => 163),
  (x => 328, y => 163),
  (x => 329, y => 163),
  (x => 330, y => 163),
  (x => 331, y => 163),
  (x => 350, y => 163),
  (x => 351, y => 163),
  (x => 352, y => 163),
  (x => 353, y => 163),
  (x => 354, y => 163),
  (x => 355, y => 163),
  (x => 356, y => 163),
  (x => 357, y => 163),
  (x => 368, y => 163),
  (x => 369, y => 163),
  (x => 370, y => 163),
  (x => 371, y => 163),
  (x => 372, y => 163),
  (x => 373, y => 163),
  (x => 378, y => 163),
  (x => 379, y => 163),
  (x => 380, y => 163),
  (x => 381, y => 163),
  (x => 382, y => 163),
  (x => 383, y => 163),
  (x => 394, y => 163),
  (x => 395, y => 163),
  (x => 396, y => 163),
  (x => 397, y => 163),
  (x => 398, y => 163),
  (x => 399, y => 163),
  (x => 424, y => 163),
  (x => 425, y => 163),
  (x => 426, y => 163),
  (x => 427, y => 163),
  (x => 428, y => 163),
  (x => 429, y => 163),
  (x => 430, y => 163),
  (x => 163, y => 164),
  (x => 164, y => 164),
  (x => 165, y => 164),
  (x => 166, y => 164),
  (x => 167, y => 164),
  (x => 168, y => 164),
  (x => 169, y => 164),
  (x => 170, y => 164),
  (x => 171, y => 164),
  (x => 187, y => 164),
  (x => 188, y => 164),
  (x => 189, y => 164),
  (x => 190, y => 164),
  (x => 191, y => 164),
  (x => 192, y => 164),
  (x => 193, y => 164),
  (x => 200, y => 164),
  (x => 201, y => 164),
  (x => 202, y => 164),
  (x => 203, y => 164),
  (x => 204, y => 164),
  (x => 205, y => 164),
  (x => 206, y => 164),
  (x => 217, y => 164),
  (x => 218, y => 164),
  (x => 219, y => 164),
  (x => 220, y => 164),
  (x => 221, y => 164),
  (x => 222, y => 164),
  (x => 231, y => 164),
  (x => 232, y => 164),
  (x => 233, y => 164),
  (x => 234, y => 164),
  (x => 235, y => 164),
  (x => 236, y => 164),
  (x => 237, y => 164),
  (x => 248, y => 164),
  (x => 249, y => 164),
  (x => 250, y => 164),
  (x => 251, y => 164),
  (x => 252, y => 164),
  (x => 253, y => 164),
  (x => 254, y => 164),
  (x => 266, y => 164),
  (x => 267, y => 164),
  (x => 268, y => 164),
  (x => 269, y => 164),
  (x => 270, y => 164),
  (x => 271, y => 164),
  (x => 272, y => 164),
  (x => 279, y => 164),
  (x => 280, y => 164),
  (x => 281, y => 164),
  (x => 282, y => 164),
  (x => 283, y => 164),
  (x => 284, y => 164),
  (x => 285, y => 164),
  (x => 325, y => 164),
  (x => 326, y => 164),
  (x => 327, y => 164),
  (x => 328, y => 164),
  (x => 329, y => 164),
  (x => 330, y => 164),
  (x => 331, y => 164),
  (x => 332, y => 164),
  (x => 349, y => 164),
  (x => 350, y => 164),
  (x => 351, y => 164),
  (x => 352, y => 164),
  (x => 353, y => 164),
  (x => 354, y => 164),
  (x => 355, y => 164),
  (x => 356, y => 164),
  (x => 368, y => 164),
  (x => 369, y => 164),
  (x => 370, y => 164),
  (x => 371, y => 164),
  (x => 372, y => 164),
  (x => 373, y => 164),
  (x => 378, y => 164),
  (x => 379, y => 164),
  (x => 380, y => 164),
  (x => 381, y => 164),
  (x => 382, y => 164),
  (x => 383, y => 164),
  (x => 394, y => 164),
  (x => 395, y => 164),
  (x => 396, y => 164),
  (x => 397, y => 164),
  (x => 398, y => 164),
  (x => 399, y => 164),
  (x => 424, y => 164),
  (x => 425, y => 164),
  (x => 426, y => 164),
  (x => 427, y => 164),
  (x => 428, y => 164),
  (x => 429, y => 164),
  (x => 430, y => 164),
  (x => 164, y => 165),
  (x => 165, y => 165),
  (x => 166, y => 165),
  (x => 167, y => 165),
  (x => 168, y => 165),
  (x => 169, y => 165),
  (x => 170, y => 165),
  (x => 171, y => 165),
  (x => 172, y => 165),
  (x => 187, y => 165),
  (x => 188, y => 165),
  (x => 189, y => 165),
  (x => 190, y => 165),
  (x => 191, y => 165),
  (x => 192, y => 165),
  (x => 193, y => 165),
  (x => 200, y => 165),
  (x => 201, y => 165),
  (x => 202, y => 165),
  (x => 203, y => 165),
  (x => 204, y => 165),
  (x => 205, y => 165),
  (x => 217, y => 165),
  (x => 218, y => 165),
  (x => 219, y => 165),
  (x => 220, y => 165),
  (x => 221, y => 165),
  (x => 222, y => 165),
  (x => 231, y => 165),
  (x => 232, y => 165),
  (x => 233, y => 165),
  (x => 234, y => 165),
  (x => 235, y => 165),
  (x => 236, y => 165),
  (x => 237, y => 165),
  (x => 248, y => 165),
  (x => 249, y => 165),
  (x => 250, y => 165),
  (x => 251, y => 165),
  (x => 252, y => 165),
  (x => 253, y => 165),
  (x => 254, y => 165),
  (x => 266, y => 165),
  (x => 267, y => 165),
  (x => 268, y => 165),
  (x => 269, y => 165),
  (x => 270, y => 165),
  (x => 271, y => 165),
  (x => 272, y => 165),
  (x => 279, y => 165),
  (x => 280, y => 165),
  (x => 281, y => 165),
  (x => 282, y => 165),
  (x => 283, y => 165),
  (x => 284, y => 165),
  (x => 285, y => 165),
  (x => 325, y => 165),
  (x => 326, y => 165),
  (x => 327, y => 165),
  (x => 328, y => 165),
  (x => 329, y => 165),
  (x => 330, y => 165),
  (x => 331, y => 165),
  (x => 332, y => 165),
  (x => 349, y => 165),
  (x => 350, y => 165),
  (x => 351, y => 165),
  (x => 352, y => 165),
  (x => 353, y => 165),
  (x => 354, y => 165),
  (x => 355, y => 165),
  (x => 356, y => 165),
  (x => 369, y => 165),
  (x => 370, y => 165),
  (x => 371, y => 165),
  (x => 372, y => 165),
  (x => 373, y => 165),
  (x => 374, y => 165),
  (x => 378, y => 165),
  (x => 379, y => 165),
  (x => 380, y => 165),
  (x => 381, y => 165),
  (x => 382, y => 165),
  (x => 383, y => 165),
  (x => 394, y => 165),
  (x => 395, y => 165),
  (x => 396, y => 165),
  (x => 397, y => 165),
  (x => 398, y => 165),
  (x => 399, y => 165),
  (x => 424, y => 165),
  (x => 425, y => 165),
  (x => 426, y => 165),
  (x => 427, y => 165),
  (x => 428, y => 165),
  (x => 429, y => 165),
  (x => 430, y => 165),
  (x => 164, y => 166),
  (x => 165, y => 166),
  (x => 166, y => 166),
  (x => 167, y => 166),
  (x => 168, y => 166),
  (x => 169, y => 166),
  (x => 170, y => 166),
  (x => 171, y => 166),
  (x => 172, y => 166),
  (x => 187, y => 166),
  (x => 188, y => 166),
  (x => 189, y => 166),
  (x => 190, y => 166),
  (x => 191, y => 166),
  (x => 192, y => 166),
  (x => 193, y => 166),
  (x => 200, y => 166),
  (x => 201, y => 166),
  (x => 202, y => 166),
  (x => 203, y => 166),
  (x => 204, y => 166),
  (x => 205, y => 166),
  (x => 216, y => 166),
  (x => 217, y => 166),
  (x => 218, y => 166),
  (x => 219, y => 166),
  (x => 220, y => 166),
  (x => 221, y => 166),
  (x => 222, y => 166),
  (x => 231, y => 166),
  (x => 232, y => 166),
  (x => 233, y => 166),
  (x => 234, y => 166),
  (x => 235, y => 166),
  (x => 236, y => 166),
  (x => 237, y => 166),
  (x => 248, y => 166),
  (x => 249, y => 166),
  (x => 250, y => 166),
  (x => 251, y => 166),
  (x => 252, y => 166),
  (x => 253, y => 166),
  (x => 254, y => 166),
  (x => 266, y => 166),
  (x => 267, y => 166),
  (x => 268, y => 166),
  (x => 269, y => 166),
  (x => 270, y => 166),
  (x => 271, y => 166),
  (x => 272, y => 166),
  (x => 279, y => 166),
  (x => 280, y => 166),
  (x => 281, y => 166),
  (x => 282, y => 166),
  (x => 283, y => 166),
  (x => 284, y => 166),
  (x => 285, y => 166),
  (x => 325, y => 166),
  (x => 326, y => 166),
  (x => 327, y => 166),
  (x => 328, y => 166),
  (x => 329, y => 166),
  (x => 330, y => 166),
  (x => 331, y => 166),
  (x => 332, y => 166),
  (x => 333, y => 166),
  (x => 348, y => 166),
  (x => 349, y => 166),
  (x => 350, y => 166),
  (x => 351, y => 166),
  (x => 352, y => 166),
  (x => 353, y => 166),
  (x => 354, y => 166),
  (x => 355, y => 166),
  (x => 356, y => 166),
  (x => 369, y => 166),
  (x => 370, y => 166),
  (x => 371, y => 166),
  (x => 372, y => 166),
  (x => 373, y => 166),
  (x => 374, y => 166),
  (x => 378, y => 166),
  (x => 379, y => 166),
  (x => 380, y => 166),
  (x => 381, y => 166),
  (x => 382, y => 166),
  (x => 394, y => 166),
  (x => 395, y => 166),
  (x => 396, y => 166),
  (x => 397, y => 166),
  (x => 398, y => 166),
  (x => 399, y => 166),
  (x => 400, y => 166),
  (x => 424, y => 166),
  (x => 425, y => 166),
  (x => 426, y => 166),
  (x => 427, y => 166),
  (x => 428, y => 166),
  (x => 429, y => 166),
  (x => 430, y => 166),
  (x => 165, y => 167),
  (x => 166, y => 167),
  (x => 167, y => 167),
  (x => 168, y => 167),
  (x => 169, y => 167),
  (x => 170, y => 167),
  (x => 171, y => 167),
  (x => 172, y => 167),
  (x => 173, y => 167),
  (x => 187, y => 167),
  (x => 188, y => 167),
  (x => 189, y => 167),
  (x => 190, y => 167),
  (x => 191, y => 167),
  (x => 192, y => 167),
  (x => 193, y => 167),
  (x => 200, y => 167),
  (x => 201, y => 167),
  (x => 202, y => 167),
  (x => 203, y => 167),
  (x => 204, y => 167),
  (x => 205, y => 167),
  (x => 216, y => 167),
  (x => 217, y => 167),
  (x => 218, y => 167),
  (x => 219, y => 167),
  (x => 220, y => 167),
  (x => 221, y => 167),
  (x => 222, y => 167),
  (x => 231, y => 167),
  (x => 232, y => 167),
  (x => 233, y => 167),
  (x => 234, y => 167),
  (x => 235, y => 167),
  (x => 236, y => 167),
  (x => 237, y => 167),
  (x => 248, y => 167),
  (x => 249, y => 167),
  (x => 250, y => 167),
  (x => 251, y => 167),
  (x => 252, y => 167),
  (x => 253, y => 167),
  (x => 254, y => 167),
  (x => 266, y => 167),
  (x => 267, y => 167),
  (x => 268, y => 167),
  (x => 269, y => 167),
  (x => 270, y => 167),
  (x => 271, y => 167),
  (x => 272, y => 167),
  (x => 280, y => 167),
  (x => 281, y => 167),
  (x => 282, y => 167),
  (x => 283, y => 167),
  (x => 284, y => 167),
  (x => 285, y => 167),
  (x => 326, y => 167),
  (x => 327, y => 167),
  (x => 328, y => 167),
  (x => 329, y => 167),
  (x => 330, y => 167),
  (x => 331, y => 167),
  (x => 332, y => 167),
  (x => 333, y => 167),
  (x => 334, y => 167),
  (x => 347, y => 167),
  (x => 348, y => 167),
  (x => 349, y => 167),
  (x => 350, y => 167),
  (x => 351, y => 167),
  (x => 352, y => 167),
  (x => 353, y => 167),
  (x => 354, y => 167),
  (x => 355, y => 167),
  (x => 369, y => 167),
  (x => 370, y => 167),
  (x => 371, y => 167),
  (x => 372, y => 167),
  (x => 373, y => 167),
  (x => 374, y => 167),
  (x => 377, y => 167),
  (x => 378, y => 167),
  (x => 379, y => 167),
  (x => 380, y => 167),
  (x => 381, y => 167),
  (x => 382, y => 167),
  (x => 394, y => 167),
  (x => 395, y => 167),
  (x => 396, y => 167),
  (x => 397, y => 167),
  (x => 398, y => 167),
  (x => 399, y => 167),
  (x => 400, y => 167),
  (x => 424, y => 167),
  (x => 425, y => 167),
  (x => 426, y => 167),
  (x => 427, y => 167),
  (x => 428, y => 167),
  (x => 429, y => 167),
  (x => 430, y => 167),
  (x => 165, y => 168),
  (x => 166, y => 168),
  (x => 167, y => 168),
  (x => 168, y => 168),
  (x => 169, y => 168),
  (x => 170, y => 168),
  (x => 171, y => 168),
  (x => 172, y => 168),
  (x => 173, y => 168),
  (x => 174, y => 168),
  (x => 187, y => 168),
  (x => 188, y => 168),
  (x => 189, y => 168),
  (x => 190, y => 168),
  (x => 191, y => 168),
  (x => 192, y => 168),
  (x => 193, y => 168),
  (x => 200, y => 168),
  (x => 201, y => 168),
  (x => 202, y => 168),
  (x => 203, y => 168),
  (x => 204, y => 168),
  (x => 205, y => 168),
  (x => 216, y => 168),
  (x => 217, y => 168),
  (x => 218, y => 168),
  (x => 219, y => 168),
  (x => 220, y => 168),
  (x => 221, y => 168),
  (x => 222, y => 168),
  (x => 231, y => 168),
  (x => 232, y => 168),
  (x => 233, y => 168),
  (x => 234, y => 168),
  (x => 235, y => 168),
  (x => 236, y => 168),
  (x => 237, y => 168),
  (x => 248, y => 168),
  (x => 249, y => 168),
  (x => 250, y => 168),
  (x => 251, y => 168),
  (x => 252, y => 168),
  (x => 253, y => 168),
  (x => 254, y => 168),
  (x => 266, y => 168),
  (x => 267, y => 168),
  (x => 268, y => 168),
  (x => 269, y => 168),
  (x => 270, y => 168),
  (x => 271, y => 168),
  (x => 272, y => 168),
  (x => 280, y => 168),
  (x => 281, y => 168),
  (x => 282, y => 168),
  (x => 283, y => 168),
  (x => 284, y => 168),
  (x => 285, y => 168),
  (x => 286, y => 168),
  (x => 326, y => 168),
  (x => 327, y => 168),
  (x => 328, y => 168),
  (x => 329, y => 168),
  (x => 330, y => 168),
  (x => 331, y => 168),
  (x => 332, y => 168),
  (x => 333, y => 168),
  (x => 334, y => 168),
  (x => 335, y => 168),
  (x => 346, y => 168),
  (x => 347, y => 168),
  (x => 348, y => 168),
  (x => 349, y => 168),
  (x => 350, y => 168),
  (x => 351, y => 168),
  (x => 352, y => 168),
  (x => 353, y => 168),
  (x => 354, y => 168),
  (x => 355, y => 168),
  (x => 369, y => 168),
  (x => 370, y => 168),
  (x => 371, y => 168),
  (x => 372, y => 168),
  (x => 373, y => 168),
  (x => 374, y => 168),
  (x => 377, y => 168),
  (x => 378, y => 168),
  (x => 379, y => 168),
  (x => 380, y => 168),
  (x => 381, y => 168),
  (x => 382, y => 168),
  (x => 394, y => 168),
  (x => 395, y => 168),
  (x => 396, y => 168),
  (x => 397, y => 168),
  (x => 398, y => 168),
  (x => 399, y => 168),
  (x => 400, y => 168),
  (x => 424, y => 168),
  (x => 425, y => 168),
  (x => 426, y => 168),
  (x => 427, y => 168),
  (x => 428, y => 168),
  (x => 429, y => 168),
  (x => 430, y => 168),
  (x => 165, y => 169),
  (x => 166, y => 169),
  (x => 167, y => 169),
  (x => 168, y => 169),
  (x => 169, y => 169),
  (x => 170, y => 169),
  (x => 171, y => 169),
  (x => 172, y => 169),
  (x => 173, y => 169),
  (x => 174, y => 169),
  (x => 175, y => 169),
  (x => 176, y => 169),
  (x => 187, y => 169),
  (x => 188, y => 169),
  (x => 189, y => 169),
  (x => 190, y => 169),
  (x => 191, y => 169),
  (x => 192, y => 169),
  (x => 193, y => 169),
  (x => 200, y => 169),
  (x => 201, y => 169),
  (x => 202, y => 169),
  (x => 203, y => 169),
  (x => 204, y => 169),
  (x => 205, y => 169),
  (x => 206, y => 169),
  (x => 215, y => 169),
  (x => 216, y => 169),
  (x => 217, y => 169),
  (x => 218, y => 169),
  (x => 219, y => 169),
  (x => 220, y => 169),
  (x => 221, y => 169),
  (x => 222, y => 169),
  (x => 231, y => 169),
  (x => 232, y => 169),
  (x => 233, y => 169),
  (x => 234, y => 169),
  (x => 235, y => 169),
  (x => 236, y => 169),
  (x => 237, y => 169),
  (x => 248, y => 169),
  (x => 249, y => 169),
  (x => 250, y => 169),
  (x => 251, y => 169),
  (x => 252, y => 169),
  (x => 253, y => 169),
  (x => 254, y => 169),
  (x => 266, y => 169),
  (x => 267, y => 169),
  (x => 268, y => 169),
  (x => 269, y => 169),
  (x => 270, y => 169),
  (x => 271, y => 169),
  (x => 272, y => 169),
  (x => 280, y => 169),
  (x => 281, y => 169),
  (x => 282, y => 169),
  (x => 283, y => 169),
  (x => 284, y => 169),
  (x => 285, y => 169),
  (x => 286, y => 169),
  (x => 327, y => 169),
  (x => 328, y => 169),
  (x => 329, y => 169),
  (x => 330, y => 169),
  (x => 331, y => 169),
  (x => 332, y => 169),
  (x => 333, y => 169),
  (x => 334, y => 169),
  (x => 335, y => 169),
  (x => 336, y => 169),
  (x => 345, y => 169),
  (x => 346, y => 169),
  (x => 347, y => 169),
  (x => 348, y => 169),
  (x => 349, y => 169),
  (x => 350, y => 169),
  (x => 351, y => 169),
  (x => 352, y => 169),
  (x => 353, y => 169),
  (x => 354, y => 169),
  (x => 370, y => 169),
  (x => 371, y => 169),
  (x => 372, y => 169),
  (x => 373, y => 169),
  (x => 374, y => 169),
  (x => 377, y => 169),
  (x => 378, y => 169),
  (x => 379, y => 169),
  (x => 380, y => 169),
  (x => 381, y => 169),
  (x => 395, y => 169),
  (x => 396, y => 169),
  (x => 397, y => 169),
  (x => 398, y => 169),
  (x => 399, y => 169),
  (x => 400, y => 169),
  (x => 401, y => 169),
  (x => 424, y => 169),
  (x => 425, y => 169),
  (x => 426, y => 169),
  (x => 427, y => 169),
  (x => 428, y => 169),
  (x => 429, y => 169),
  (x => 430, y => 169),
  (x => 166, y => 170),
  (x => 167, y => 170),
  (x => 168, y => 170),
  (x => 169, y => 170),
  (x => 170, y => 170),
  (x => 171, y => 170),
  (x => 172, y => 170),
  (x => 173, y => 170),
  (x => 174, y => 170),
  (x => 175, y => 170),
  (x => 176, y => 170),
  (x => 177, y => 170),
  (x => 178, y => 170),
  (x => 184, y => 170),
  (x => 185, y => 170),
  (x => 186, y => 170),
  (x => 187, y => 170),
  (x => 188, y => 170),
  (x => 189, y => 170),
  (x => 190, y => 170),
  (x => 191, y => 170),
  (x => 192, y => 170),
  (x => 193, y => 170),
  (x => 200, y => 170),
  (x => 201, y => 170),
  (x => 202, y => 170),
  (x => 203, y => 170),
  (x => 204, y => 170),
  (x => 205, y => 170),
  (x => 206, y => 170),
  (x => 214, y => 170),
  (x => 215, y => 170),
  (x => 216, y => 170),
  (x => 217, y => 170),
  (x => 218, y => 170),
  (x => 219, y => 170),
  (x => 220, y => 170),
  (x => 221, y => 170),
  (x => 222, y => 170),
  (x => 231, y => 170),
  (x => 232, y => 170),
  (x => 233, y => 170),
  (x => 234, y => 170),
  (x => 235, y => 170),
  (x => 236, y => 170),
  (x => 237, y => 170),
  (x => 248, y => 170),
  (x => 249, y => 170),
  (x => 250, y => 170),
  (x => 251, y => 170),
  (x => 252, y => 170),
  (x => 253, y => 170),
  (x => 254, y => 170),
  (x => 266, y => 170),
  (x => 267, y => 170),
  (x => 268, y => 170),
  (x => 269, y => 170),
  (x => 270, y => 170),
  (x => 271, y => 170),
  (x => 272, y => 170),
  (x => 280, y => 170),
  (x => 281, y => 170),
  (x => 282, y => 170),
  (x => 283, y => 170),
  (x => 284, y => 170),
  (x => 285, y => 170),
  (x => 286, y => 170),
  (x => 287, y => 170),
  (x => 327, y => 170),
  (x => 328, y => 170),
  (x => 329, y => 170),
  (x => 330, y => 170),
  (x => 331, y => 170),
  (x => 332, y => 170),
  (x => 333, y => 170),
  (x => 334, y => 170),
  (x => 335, y => 170),
  (x => 336, y => 170),
  (x => 337, y => 170),
  (x => 338, y => 170),
  (x => 339, y => 170),
  (x => 340, y => 170),
  (x => 341, y => 170),
  (x => 342, y => 170),
  (x => 343, y => 170),
  (x => 344, y => 170),
  (x => 345, y => 170),
  (x => 346, y => 170),
  (x => 347, y => 170),
  (x => 348, y => 170),
  (x => 349, y => 170),
  (x => 350, y => 170),
  (x => 351, y => 170),
  (x => 352, y => 170),
  (x => 353, y => 170),
  (x => 354, y => 170),
  (x => 370, y => 170),
  (x => 371, y => 170),
  (x => 372, y => 170),
  (x => 373, y => 170),
  (x => 374, y => 170),
  (x => 377, y => 170),
  (x => 378, y => 170),
  (x => 379, y => 170),
  (x => 380, y => 170),
  (x => 381, y => 170),
  (x => 395, y => 170),
  (x => 396, y => 170),
  (x => 397, y => 170),
  (x => 398, y => 170),
  (x => 399, y => 170),
  (x => 400, y => 170),
  (x => 401, y => 170),
  (x => 402, y => 170),
  (x => 415, y => 170),
  (x => 424, y => 170),
  (x => 425, y => 170),
  (x => 426, y => 170),
  (x => 427, y => 170),
  (x => 428, y => 170),
  (x => 429, y => 170),
  (x => 430, y => 170),
  (x => 167, y => 171),
  (x => 168, y => 171),
  (x => 169, y => 171),
  (x => 170, y => 171),
  (x => 171, y => 171),
  (x => 172, y => 171),
  (x => 173, y => 171),
  (x => 174, y => 171),
  (x => 175, y => 171),
  (x => 176, y => 171),
  (x => 177, y => 171),
  (x => 178, y => 171),
  (x => 179, y => 171),
  (x => 180, y => 171),
  (x => 181, y => 171),
  (x => 182, y => 171),
  (x => 183, y => 171),
  (x => 184, y => 171),
  (x => 185, y => 171),
  (x => 186, y => 171),
  (x => 187, y => 171),
  (x => 188, y => 171),
  (x => 189, y => 171),
  (x => 190, y => 171),
  (x => 191, y => 171),
  (x => 192, y => 171),
  (x => 193, y => 171),
  (x => 200, y => 171),
  (x => 201, y => 171),
  (x => 202, y => 171),
  (x => 203, y => 171),
  (x => 204, y => 171),
  (x => 205, y => 171),
  (x => 206, y => 171),
  (x => 207, y => 171),
  (x => 213, y => 171),
  (x => 214, y => 171),
  (x => 215, y => 171),
  (x => 216, y => 171),
  (x => 217, y => 171),
  (x => 218, y => 171),
  (x => 219, y => 171),
  (x => 220, y => 171),
  (x => 221, y => 171),
  (x => 222, y => 171),
  (x => 231, y => 171),
  (x => 232, y => 171),
  (x => 233, y => 171),
  (x => 234, y => 171),
  (x => 235, y => 171),
  (x => 236, y => 171),
  (x => 237, y => 171),
  (x => 248, y => 171),
  (x => 249, y => 171),
  (x => 250, y => 171),
  (x => 251, y => 171),
  (x => 252, y => 171),
  (x => 253, y => 171),
  (x => 254, y => 171),
  (x => 266, y => 171),
  (x => 267, y => 171),
  (x => 268, y => 171),
  (x => 269, y => 171),
  (x => 270, y => 171),
  (x => 271, y => 171),
  (x => 272, y => 171),
  (x => 281, y => 171),
  (x => 282, y => 171),
  (x => 283, y => 171),
  (x => 284, y => 171),
  (x => 285, y => 171),
  (x => 286, y => 171),
  (x => 287, y => 171),
  (x => 288, y => 171),
  (x => 289, y => 171),
  (x => 299, y => 171),
  (x => 300, y => 171),
  (x => 328, y => 171),
  (x => 329, y => 171),
  (x => 330, y => 171),
  (x => 331, y => 171),
  (x => 332, y => 171),
  (x => 333, y => 171),
  (x => 334, y => 171),
  (x => 335, y => 171),
  (x => 336, y => 171),
  (x => 337, y => 171),
  (x => 338, y => 171),
  (x => 339, y => 171),
  (x => 340, y => 171),
  (x => 341, y => 171),
  (x => 342, y => 171),
  (x => 343, y => 171),
  (x => 344, y => 171),
  (x => 345, y => 171),
  (x => 346, y => 171),
  (x => 347, y => 171),
  (x => 348, y => 171),
  (x => 349, y => 171),
  (x => 350, y => 171),
  (x => 351, y => 171),
  (x => 352, y => 171),
  (x => 353, y => 171),
  (x => 370, y => 171),
  (x => 371, y => 171),
  (x => 372, y => 171),
  (x => 373, y => 171),
  (x => 374, y => 171),
  (x => 375, y => 171),
  (x => 376, y => 171),
  (x => 377, y => 171),
  (x => 378, y => 171),
  (x => 379, y => 171),
  (x => 380, y => 171),
  (x => 381, y => 171),
  (x => 395, y => 171),
  (x => 396, y => 171),
  (x => 397, y => 171),
  (x => 398, y => 171),
  (x => 399, y => 171),
  (x => 400, y => 171),
  (x => 401, y => 171),
  (x => 402, y => 171),
  (x => 403, y => 171),
  (x => 413, y => 171),
  (x => 414, y => 171),
  (x => 415, y => 171),
  (x => 424, y => 171),
  (x => 425, y => 171),
  (x => 426, y => 171),
  (x => 427, y => 171),
  (x => 428, y => 171),
  (x => 429, y => 171),
  (x => 430, y => 171),
  (x => 167, y => 172),
  (x => 168, y => 172),
  (x => 169, y => 172),
  (x => 170, y => 172),
  (x => 171, y => 172),
  (x => 172, y => 172),
  (x => 173, y => 172),
  (x => 174, y => 172),
  (x => 175, y => 172),
  (x => 176, y => 172),
  (x => 177, y => 172),
  (x => 178, y => 172),
  (x => 179, y => 172),
  (x => 180, y => 172),
  (x => 181, y => 172),
  (x => 182, y => 172),
  (x => 183, y => 172),
  (x => 184, y => 172),
  (x => 185, y => 172),
  (x => 186, y => 172),
  (x => 187, y => 172),
  (x => 188, y => 172),
  (x => 189, y => 172),
  (x => 190, y => 172),
  (x => 191, y => 172),
  (x => 192, y => 172),
  (x => 193, y => 172),
  (x => 200, y => 172),
  (x => 201, y => 172),
  (x => 202, y => 172),
  (x => 203, y => 172),
  (x => 204, y => 172),
  (x => 205, y => 172),
  (x => 206, y => 172),
  (x => 207, y => 172),
  (x => 208, y => 172),
  (x => 209, y => 172),
  (x => 210, y => 172),
  (x => 211, y => 172),
  (x => 212, y => 172),
  (x => 213, y => 172),
  (x => 214, y => 172),
  (x => 215, y => 172),
  (x => 216, y => 172),
  (x => 217, y => 172),
  (x => 218, y => 172),
  (x => 219, y => 172),
  (x => 220, y => 172),
  (x => 221, y => 172),
  (x => 222, y => 172),
  (x => 231, y => 172),
  (x => 232, y => 172),
  (x => 233, y => 172),
  (x => 234, y => 172),
  (x => 235, y => 172),
  (x => 236, y => 172),
  (x => 237, y => 172),
  (x => 248, y => 172),
  (x => 249, y => 172),
  (x => 250, y => 172),
  (x => 251, y => 172),
  (x => 252, y => 172),
  (x => 253, y => 172),
  (x => 254, y => 172),
  (x => 266, y => 172),
  (x => 267, y => 172),
  (x => 268, y => 172),
  (x => 269, y => 172),
  (x => 270, y => 172),
  (x => 271, y => 172),
  (x => 272, y => 172),
  (x => 281, y => 172),
  (x => 282, y => 172),
  (x => 283, y => 172),
  (x => 284, y => 172),
  (x => 285, y => 172),
  (x => 286, y => 172),
  (x => 287, y => 172),
  (x => 288, y => 172),
  (x => 289, y => 172),
  (x => 290, y => 172),
  (x => 291, y => 172),
  (x => 292, y => 172),
  (x => 293, y => 172),
  (x => 294, y => 172),
  (x => 295, y => 172),
  (x => 296, y => 172),
  (x => 297, y => 172),
  (x => 298, y => 172),
  (x => 299, y => 172),
  (x => 300, y => 172),
  (x => 329, y => 172),
  (x => 330, y => 172),
  (x => 331, y => 172),
  (x => 332, y => 172),
  (x => 333, y => 172),
  (x => 334, y => 172),
  (x => 335, y => 172),
  (x => 336, y => 172),
  (x => 337, y => 172),
  (x => 338, y => 172),
  (x => 339, y => 172),
  (x => 340, y => 172),
  (x => 341, y => 172),
  (x => 342, y => 172),
  (x => 343, y => 172),
  (x => 344, y => 172),
  (x => 345, y => 172),
  (x => 346, y => 172),
  (x => 347, y => 172),
  (x => 348, y => 172),
  (x => 349, y => 172),
  (x => 350, y => 172),
  (x => 351, y => 172),
  (x => 352, y => 172),
  (x => 370, y => 172),
  (x => 371, y => 172),
  (x => 372, y => 172),
  (x => 373, y => 172),
  (x => 374, y => 172),
  (x => 375, y => 172),
  (x => 376, y => 172),
  (x => 377, y => 172),
  (x => 378, y => 172),
  (x => 379, y => 172),
  (x => 380, y => 172),
  (x => 381, y => 172),
  (x => 396, y => 172),
  (x => 397, y => 172),
  (x => 398, y => 172),
  (x => 399, y => 172),
  (x => 400, y => 172),
  (x => 401, y => 172),
  (x => 402, y => 172),
  (x => 403, y => 172),
  (x => 404, y => 172),
  (x => 405, y => 172),
  (x => 406, y => 172),
  (x => 407, y => 172),
  (x => 408, y => 172),
  (x => 409, y => 172),
  (x => 410, y => 172),
  (x => 411, y => 172),
  (x => 412, y => 172),
  (x => 413, y => 172),
  (x => 414, y => 172),
  (x => 415, y => 172),
  (x => 424, y => 172),
  (x => 425, y => 172),
  (x => 426, y => 172),
  (x => 427, y => 172),
  (x => 428, y => 172),
  (x => 429, y => 172),
  (x => 430, y => 172),
  (x => 168, y => 173),
  (x => 169, y => 173),
  (x => 170, y => 173),
  (x => 171, y => 173),
  (x => 172, y => 173),
  (x => 173, y => 173),
  (x => 174, y => 173),
  (x => 175, y => 173),
  (x => 176, y => 173),
  (x => 177, y => 173),
  (x => 178, y => 173),
  (x => 179, y => 173),
  (x => 180, y => 173),
  (x => 181, y => 173),
  (x => 182, y => 173),
  (x => 183, y => 173),
  (x => 184, y => 173),
  (x => 185, y => 173),
  (x => 186, y => 173),
  (x => 187, y => 173),
  (x => 188, y => 173),
  (x => 189, y => 173),
  (x => 190, y => 173),
  (x => 191, y => 173),
  (x => 192, y => 173),
  (x => 193, y => 173),
  (x => 201, y => 173),
  (x => 202, y => 173),
  (x => 203, y => 173),
  (x => 204, y => 173),
  (x => 205, y => 173),
  (x => 206, y => 173),
  (x => 207, y => 173),
  (x => 208, y => 173),
  (x => 209, y => 173),
  (x => 210, y => 173),
  (x => 211, y => 173),
  (x => 212, y => 173),
  (x => 213, y => 173),
  (x => 214, y => 173),
  (x => 217, y => 173),
  (x => 218, y => 173),
  (x => 219, y => 173),
  (x => 220, y => 173),
  (x => 221, y => 173),
  (x => 222, y => 173),
  (x => 231, y => 173),
  (x => 232, y => 173),
  (x => 233, y => 173),
  (x => 234, y => 173),
  (x => 235, y => 173),
  (x => 236, y => 173),
  (x => 237, y => 173),
  (x => 248, y => 173),
  (x => 249, y => 173),
  (x => 250, y => 173),
  (x => 251, y => 173),
  (x => 252, y => 173),
  (x => 253, y => 173),
  (x => 254, y => 173),
  (x => 266, y => 173),
  (x => 267, y => 173),
  (x => 268, y => 173),
  (x => 269, y => 173),
  (x => 270, y => 173),
  (x => 271, y => 173),
  (x => 272, y => 173),
  (x => 282, y => 173),
  (x => 283, y => 173),
  (x => 284, y => 173),
  (x => 285, y => 173),
  (x => 286, y => 173),
  (x => 287, y => 173),
  (x => 288, y => 173),
  (x => 289, y => 173),
  (x => 290, y => 173),
  (x => 291, y => 173),
  (x => 292, y => 173),
  (x => 293, y => 173),
  (x => 294, y => 173),
  (x => 295, y => 173),
  (x => 296, y => 173),
  (x => 297, y => 173),
  (x => 298, y => 173),
  (x => 299, y => 173),
  (x => 300, y => 173),
  (x => 329, y => 173),
  (x => 330, y => 173),
  (x => 331, y => 173),
  (x => 332, y => 173),
  (x => 333, y => 173),
  (x => 334, y => 173),
  (x => 335, y => 173),
  (x => 336, y => 173),
  (x => 337, y => 173),
  (x => 338, y => 173),
  (x => 339, y => 173),
  (x => 340, y => 173),
  (x => 341, y => 173),
  (x => 342, y => 173),
  (x => 343, y => 173),
  (x => 344, y => 173),
  (x => 345, y => 173),
  (x => 346, y => 173),
  (x => 347, y => 173),
  (x => 348, y => 173),
  (x => 349, y => 173),
  (x => 350, y => 173),
  (x => 351, y => 173),
  (x => 371, y => 173),
  (x => 372, y => 173),
  (x => 373, y => 173),
  (x => 374, y => 173),
  (x => 375, y => 173),
  (x => 376, y => 173),
  (x => 377, y => 173),
  (x => 378, y => 173),
  (x => 379, y => 173),
  (x => 380, y => 173),
  (x => 396, y => 173),
  (x => 397, y => 173),
  (x => 398, y => 173),
  (x => 399, y => 173),
  (x => 400, y => 173),
  (x => 401, y => 173),
  (x => 402, y => 173),
  (x => 403, y => 173),
  (x => 404, y => 173),
  (x => 405, y => 173),
  (x => 406, y => 173),
  (x => 407, y => 173),
  (x => 408, y => 173),
  (x => 409, y => 173),
  (x => 410, y => 173),
  (x => 411, y => 173),
  (x => 412, y => 173),
  (x => 413, y => 173),
  (x => 414, y => 173),
  (x => 415, y => 173),
  (x => 424, y => 173),
  (x => 425, y => 173),
  (x => 426, y => 173),
  (x => 427, y => 173),
  (x => 428, y => 173),
  (x => 429, y => 173),
  (x => 430, y => 173),
  (x => 169, y => 174),
  (x => 170, y => 174),
  (x => 171, y => 174),
  (x => 172, y => 174),
  (x => 173, y => 174),
  (x => 174, y => 174),
  (x => 175, y => 174),
  (x => 176, y => 174),
  (x => 177, y => 174),
  (x => 178, y => 174),
  (x => 179, y => 174),
  (x => 180, y => 174),
  (x => 181, y => 174),
  (x => 182, y => 174),
  (x => 183, y => 174),
  (x => 184, y => 174),
  (x => 185, y => 174),
  (x => 186, y => 174),
  (x => 187, y => 174),
  (x => 188, y => 174),
  (x => 189, y => 174),
  (x => 190, y => 174),
  (x => 191, y => 174),
  (x => 192, y => 174),
  (x => 193, y => 174),
  (x => 201, y => 174),
  (x => 202, y => 174),
  (x => 203, y => 174),
  (x => 204, y => 174),
  (x => 205, y => 174),
  (x => 206, y => 174),
  (x => 207, y => 174),
  (x => 208, y => 174),
  (x => 209, y => 174),
  (x => 210, y => 174),
  (x => 211, y => 174),
  (x => 212, y => 174),
  (x => 213, y => 174),
  (x => 217, y => 174),
  (x => 218, y => 174),
  (x => 219, y => 174),
  (x => 220, y => 174),
  (x => 221, y => 174),
  (x => 222, y => 174),
  (x => 231, y => 174),
  (x => 232, y => 174),
  (x => 233, y => 174),
  (x => 234, y => 174),
  (x => 235, y => 174),
  (x => 236, y => 174),
  (x => 237, y => 174),
  (x => 248, y => 174),
  (x => 249, y => 174),
  (x => 250, y => 174),
  (x => 251, y => 174),
  (x => 252, y => 174),
  (x => 253, y => 174),
  (x => 254, y => 174),
  (x => 266, y => 174),
  (x => 267, y => 174),
  (x => 268, y => 174),
  (x => 269, y => 174),
  (x => 270, y => 174),
  (x => 271, y => 174),
  (x => 272, y => 174),
  (x => 283, y => 174),
  (x => 284, y => 174),
  (x => 285, y => 174),
  (x => 286, y => 174),
  (x => 287, y => 174),
  (x => 288, y => 174),
  (x => 289, y => 174),
  (x => 290, y => 174),
  (x => 291, y => 174),
  (x => 292, y => 174),
  (x => 293, y => 174),
  (x => 294, y => 174),
  (x => 295, y => 174),
  (x => 296, y => 174),
  (x => 297, y => 174),
  (x => 298, y => 174),
  (x => 299, y => 174),
  (x => 300, y => 174),
  (x => 330, y => 174),
  (x => 331, y => 174),
  (x => 332, y => 174),
  (x => 333, y => 174),
  (x => 334, y => 174),
  (x => 335, y => 174),
  (x => 336, y => 174),
  (x => 337, y => 174),
  (x => 338, y => 174),
  (x => 339, y => 174),
  (x => 340, y => 174),
  (x => 341, y => 174),
  (x => 342, y => 174),
  (x => 343, y => 174),
  (x => 344, y => 174),
  (x => 345, y => 174),
  (x => 346, y => 174),
  (x => 347, y => 174),
  (x => 348, y => 174),
  (x => 349, y => 174),
  (x => 350, y => 174),
  (x => 351, y => 174),
  (x => 371, y => 174),
  (x => 372, y => 174),
  (x => 373, y => 174),
  (x => 374, y => 174),
  (x => 375, y => 174),
  (x => 376, y => 174),
  (x => 377, y => 174),
  (x => 378, y => 174),
  (x => 379, y => 174),
  (x => 380, y => 174),
  (x => 397, y => 174),
  (x => 398, y => 174),
  (x => 399, y => 174),
  (x => 400, y => 174),
  (x => 401, y => 174),
  (x => 402, y => 174),
  (x => 403, y => 174),
  (x => 404, y => 174),
  (x => 405, y => 174),
  (x => 406, y => 174),
  (x => 407, y => 174),
  (x => 408, y => 174),
  (x => 409, y => 174),
  (x => 410, y => 174),
  (x => 411, y => 174),
  (x => 412, y => 174),
  (x => 413, y => 174),
  (x => 414, y => 174),
  (x => 415, y => 174),
  (x => 424, y => 174),
  (x => 425, y => 174),
  (x => 426, y => 174),
  (x => 427, y => 174),
  (x => 428, y => 174),
  (x => 429, y => 174),
  (x => 430, y => 174),
  (x => 171, y => 175),
  (x => 172, y => 175),
  (x => 173, y => 175),
  (x => 174, y => 175),
  (x => 175, y => 175),
  (x => 176, y => 175),
  (x => 177, y => 175),
  (x => 178, y => 175),
  (x => 179, y => 175),
  (x => 180, y => 175),
  (x => 181, y => 175),
  (x => 182, y => 175),
  (x => 183, y => 175),
  (x => 184, y => 175),
  (x => 185, y => 175),
  (x => 186, y => 175),
  (x => 187, y => 175),
  (x => 188, y => 175),
  (x => 189, y => 175),
  (x => 190, y => 175),
  (x => 191, y => 175),
  (x => 192, y => 175),
  (x => 202, y => 175),
  (x => 203, y => 175),
  (x => 204, y => 175),
  (x => 205, y => 175),
  (x => 206, y => 175),
  (x => 207, y => 175),
  (x => 208, y => 175),
  (x => 209, y => 175),
  (x => 210, y => 175),
  (x => 211, y => 175),
  (x => 212, y => 175),
  (x => 213, y => 175),
  (x => 217, y => 175),
  (x => 218, y => 175),
  (x => 219, y => 175),
  (x => 220, y => 175),
  (x => 221, y => 175),
  (x => 222, y => 175),
  (x => 231, y => 175),
  (x => 232, y => 175),
  (x => 233, y => 175),
  (x => 234, y => 175),
  (x => 235, y => 175),
  (x => 236, y => 175),
  (x => 237, y => 175),
  (x => 248, y => 175),
  (x => 249, y => 175),
  (x => 250, y => 175),
  (x => 251, y => 175),
  (x => 252, y => 175),
  (x => 253, y => 175),
  (x => 254, y => 175),
  (x => 266, y => 175),
  (x => 267, y => 175),
  (x => 268, y => 175),
  (x => 269, y => 175),
  (x => 270, y => 175),
  (x => 271, y => 175),
  (x => 272, y => 175),
  (x => 283, y => 175),
  (x => 284, y => 175),
  (x => 285, y => 175),
  (x => 286, y => 175),
  (x => 287, y => 175),
  (x => 288, y => 175),
  (x => 289, y => 175),
  (x => 290, y => 175),
  (x => 291, y => 175),
  (x => 292, y => 175),
  (x => 293, y => 175),
  (x => 294, y => 175),
  (x => 295, y => 175),
  (x => 296, y => 175),
  (x => 297, y => 175),
  (x => 298, y => 175),
  (x => 299, y => 175),
  (x => 300, y => 175),
  (x => 331, y => 175),
  (x => 332, y => 175),
  (x => 333, y => 175),
  (x => 334, y => 175),
  (x => 335, y => 175),
  (x => 336, y => 175),
  (x => 337, y => 175),
  (x => 338, y => 175),
  (x => 339, y => 175),
  (x => 340, y => 175),
  (x => 341, y => 175),
  (x => 342, y => 175),
  (x => 343, y => 175),
  (x => 344, y => 175),
  (x => 345, y => 175),
  (x => 346, y => 175),
  (x => 347, y => 175),
  (x => 348, y => 175),
  (x => 349, y => 175),
  (x => 371, y => 175),
  (x => 372, y => 175),
  (x => 373, y => 175),
  (x => 374, y => 175),
  (x => 375, y => 175),
  (x => 376, y => 175),
  (x => 377, y => 175),
  (x => 378, y => 175),
  (x => 379, y => 175),
  (x => 380, y => 175),
  (x => 398, y => 175),
  (x => 399, y => 175),
  (x => 400, y => 175),
  (x => 401, y => 175),
  (x => 402, y => 175),
  (x => 403, y => 175),
  (x => 404, y => 175),
  (x => 405, y => 175),
  (x => 406, y => 175),
  (x => 407, y => 175),
  (x => 408, y => 175),
  (x => 409, y => 175),
  (x => 410, y => 175),
  (x => 411, y => 175),
  (x => 412, y => 175),
  (x => 413, y => 175),
  (x => 414, y => 175),
  (x => 415, y => 175),
  (x => 424, y => 175),
  (x => 425, y => 175),
  (x => 426, y => 175),
  (x => 427, y => 175),
  (x => 428, y => 175),
  (x => 429, y => 175),
  (x => 430, y => 175),
  (x => 172, y => 176),
  (x => 173, y => 176),
  (x => 174, y => 176),
  (x => 175, y => 176),
  (x => 176, y => 176),
  (x => 177, y => 176),
  (x => 178, y => 176),
  (x => 179, y => 176),
  (x => 180, y => 176),
  (x => 181, y => 176),
  (x => 182, y => 176),
  (x => 183, y => 176),
  (x => 184, y => 176),
  (x => 185, y => 176),
  (x => 186, y => 176),
  (x => 187, y => 176),
  (x => 188, y => 176),
  (x => 189, y => 176),
  (x => 190, y => 176),
  (x => 202, y => 176),
  (x => 203, y => 176),
  (x => 204, y => 176),
  (x => 205, y => 176),
  (x => 206, y => 176),
  (x => 207, y => 176),
  (x => 208, y => 176),
  (x => 209, y => 176),
  (x => 210, y => 176),
  (x => 211, y => 176),
  (x => 212, y => 176),
  (x => 217, y => 176),
  (x => 218, y => 176),
  (x => 219, y => 176),
  (x => 220, y => 176),
  (x => 221, y => 176),
  (x => 222, y => 176),
  (x => 231, y => 176),
  (x => 232, y => 176),
  (x => 233, y => 176),
  (x => 234, y => 176),
  (x => 235, y => 176),
  (x => 236, y => 176),
  (x => 237, y => 176),
  (x => 248, y => 176),
  (x => 249, y => 176),
  (x => 250, y => 176),
  (x => 251, y => 176),
  (x => 252, y => 176),
  (x => 253, y => 176),
  (x => 254, y => 176),
  (x => 266, y => 176),
  (x => 267, y => 176),
  (x => 268, y => 176),
  (x => 269, y => 176),
  (x => 270, y => 176),
  (x => 271, y => 176),
  (x => 272, y => 176),
  (x => 285, y => 176),
  (x => 286, y => 176),
  (x => 287, y => 176),
  (x => 288, y => 176),
  (x => 289, y => 176),
  (x => 290, y => 176),
  (x => 291, y => 176),
  (x => 292, y => 176),
  (x => 293, y => 176),
  (x => 294, y => 176),
  (x => 295, y => 176),
  (x => 296, y => 176),
  (x => 297, y => 176),
  (x => 298, y => 176),
  (x => 299, y => 176),
  (x => 300, y => 176),
  (x => 333, y => 176),
  (x => 334, y => 176),
  (x => 335, y => 176),
  (x => 336, y => 176),
  (x => 337, y => 176),
  (x => 338, y => 176),
  (x => 339, y => 176),
  (x => 340, y => 176),
  (x => 341, y => 176),
  (x => 342, y => 176),
  (x => 343, y => 176),
  (x => 344, y => 176),
  (x => 345, y => 176),
  (x => 346, y => 176),
  (x => 347, y => 176),
  (x => 348, y => 176),
  (x => 371, y => 176),
  (x => 372, y => 176),
  (x => 373, y => 176),
  (x => 374, y => 176),
  (x => 375, y => 176),
  (x => 376, y => 176),
  (x => 377, y => 176),
  (x => 378, y => 176),
  (x => 379, y => 176),
  (x => 399, y => 176),
  (x => 400, y => 176),
  (x => 401, y => 176),
  (x => 402, y => 176),
  (x => 403, y => 176),
  (x => 404, y => 176),
  (x => 405, y => 176),
  (x => 406, y => 176),
  (x => 407, y => 176),
  (x => 408, y => 176),
  (x => 409, y => 176),
  (x => 410, y => 176),
  (x => 411, y => 176),
  (x => 412, y => 176),
  (x => 413, y => 176),
  (x => 414, y => 176),
  (x => 424, y => 176),
  (x => 425, y => 176),
  (x => 426, y => 176),
  (x => 427, y => 176),
  (x => 428, y => 176),
  (x => 429, y => 176),
  (x => 430, y => 176),
  (x => 174, y => 177),
  (x => 175, y => 177),
  (x => 176, y => 177),
  (x => 177, y => 177),
  (x => 178, y => 177),
  (x => 179, y => 177),
  (x => 180, y => 177),
  (x => 181, y => 177),
  (x => 182, y => 177),
  (x => 183, y => 177),
  (x => 184, y => 177),
  (x => 185, y => 177),
  (x => 186, y => 177),
  (x => 187, y => 177),
  (x => 188, y => 177),
  (x => 204, y => 177),
  (x => 205, y => 177),
  (x => 206, y => 177),
  (x => 207, y => 177),
  (x => 208, y => 177),
  (x => 209, y => 177),
  (x => 210, y => 177),
  (x => 211, y => 177),
  (x => 216, y => 177),
  (x => 217, y => 177),
  (x => 218, y => 177),
  (x => 219, y => 177),
  (x => 220, y => 177),
  (x => 221, y => 177),
  (x => 222, y => 177),
  (x => 231, y => 177),
  (x => 232, y => 177),
  (x => 233, y => 177),
  (x => 234, y => 177),
  (x => 235, y => 177),
  (x => 236, y => 177),
  (x => 237, y => 177),
  (x => 248, y => 177),
  (x => 249, y => 177),
  (x => 250, y => 177),
  (x => 251, y => 177),
  (x => 252, y => 177),
  (x => 253, y => 177),
  (x => 254, y => 177),
  (x => 265, y => 177),
  (x => 266, y => 177),
  (x => 267, y => 177),
  (x => 268, y => 177),
  (x => 269, y => 177),
  (x => 270, y => 177),
  (x => 271, y => 177),
  (x => 272, y => 177),
  (x => 286, y => 177),
  (x => 287, y => 177),
  (x => 288, y => 177),
  (x => 289, y => 177),
  (x => 290, y => 177),
  (x => 291, y => 177),
  (x => 292, y => 177),
  (x => 293, y => 177),
  (x => 294, y => 177),
  (x => 295, y => 177),
  (x => 296, y => 177),
  (x => 297, y => 177),
  (x => 298, y => 177),
  (x => 335, y => 177),
  (x => 336, y => 177),
  (x => 337, y => 177),
  (x => 338, y => 177),
  (x => 339, y => 177),
  (x => 340, y => 177),
  (x => 341, y => 177),
  (x => 342, y => 177),
  (x => 343, y => 177),
  (x => 344, y => 177),
  (x => 345, y => 177),
  (x => 346, y => 177),
  (x => 372, y => 177),
  (x => 373, y => 177),
  (x => 374, y => 177),
  (x => 375, y => 177),
  (x => 376, y => 177),
  (x => 377, y => 177),
  (x => 378, y => 177),
  (x => 379, y => 177),
  (x => 401, y => 177),
  (x => 402, y => 177),
  (x => 403, y => 177),
  (x => 404, y => 177),
  (x => 405, y => 177),
  (x => 406, y => 177),
  (x => 407, y => 177),
  (x => 408, y => 177),
  (x => 409, y => 177),
  (x => 410, y => 177),
  (x => 411, y => 177),
  (x => 412, y => 177),
  (x => 424, y => 177),
  (x => 425, y => 177),
  (x => 426, y => 177),
  (x => 427, y => 177),
  (x => 428, y => 177),
  (x => 429, y => 177),
  (x => 430, y => 177),
  (x => 178, y => 178),
  (x => 179, y => 178),
  (x => 180, y => 178),
  (x => 181, y => 178),
  (x => 182, y => 178),
  (x => 183, y => 178),
  (x => 206, y => 178),
  (x => 207, y => 178),
  (x => 208, y => 178),
  (x => 290, y => 178),
  (x => 291, y => 178),
  (x => 292, y => 178),
  (x => 293, y => 178),
  (x => 294, y => 178),
  (x => 338, y => 178),
  (x => 339, y => 178),
  (x => 340, y => 178),
  (x => 341, y => 178),
  (x => 342, y => 178),
  (x => 404, y => 178),
  (x => 405, y => 178),
  (x => 406, y => 178),
  (x => 407, y => 178),
  (x => 408, y => 178),
  (x => 409, y => 178),
  (x => 228, y => 222),
  (x => 229, y => 222),
  (x => 230, y => 222),
  (x => 231, y => 222),
  (x => 368, y => 222),
  (x => 369, y => 222),
  (x => 209, y => 223),
  (x => 210, y => 223),
  (x => 211, y => 223),
  (x => 212, y => 223),
  (x => 213, y => 223),
  (x => 214, y => 223),
  (x => 215, y => 223),
  (x => 216, y => 223),
  (x => 217, y => 223),
  (x => 228, y => 223),
  (x => 229, y => 223),
  (x => 230, y => 223),
  (x => 231, y => 223),
  (x => 316, y => 223),
  (x => 317, y => 223),
  (x => 334, y => 223),
  (x => 335, y => 223),
  (x => 336, y => 223),
  (x => 337, y => 223),
  (x => 347, y => 223),
  (x => 348, y => 223),
  (x => 349, y => 223),
  (x => 350, y => 223),
  (x => 360, y => 223),
  (x => 361, y => 223),
  (x => 362, y => 223),
  (x => 367, y => 223),
  (x => 368, y => 223),
  (x => 369, y => 223),
  (x => 370, y => 223),
  (x => 209, y => 224),
  (x => 210, y => 224),
  (x => 211, y => 224),
  (x => 212, y => 224),
  (x => 213, y => 224),
  (x => 214, y => 224),
  (x => 215, y => 224),
  (x => 216, y => 224),
  (x => 217, y => 224),
  (x => 218, y => 224),
  (x => 219, y => 224),
  (x => 220, y => 224),
  (x => 228, y => 224),
  (x => 229, y => 224),
  (x => 230, y => 224),
  (x => 231, y => 224),
  (x => 315, y => 224),
  (x => 316, y => 224),
  (x => 317, y => 224),
  (x => 334, y => 224),
  (x => 335, y => 224),
  (x => 336, y => 224),
  (x => 337, y => 224),
  (x => 347, y => 224),
  (x => 348, y => 224),
  (x => 349, y => 224),
  (x => 350, y => 224),
  (x => 360, y => 224),
  (x => 361, y => 224),
  (x => 362, y => 224),
  (x => 367, y => 224),
  (x => 368, y => 224),
  (x => 369, y => 224),
  (x => 370, y => 224),
  (x => 209, y => 225),
  (x => 210, y => 225),
  (x => 211, y => 225),
  (x => 212, y => 225),
  (x => 213, y => 225),
  (x => 214, y => 225),
  (x => 215, y => 225),
  (x => 216, y => 225),
  (x => 217, y => 225),
  (x => 218, y => 225),
  (x => 219, y => 225),
  (x => 220, y => 225),
  (x => 221, y => 225),
  (x => 228, y => 225),
  (x => 229, y => 225),
  (x => 230, y => 225),
  (x => 231, y => 225),
  (x => 313, y => 225),
  (x => 314, y => 225),
  (x => 315, y => 225),
  (x => 316, y => 225),
  (x => 317, y => 225),
  (x => 335, y => 225),
  (x => 336, y => 225),
  (x => 337, y => 225),
  (x => 347, y => 225),
  (x => 348, y => 225),
  (x => 349, y => 225),
  (x => 350, y => 225),
  (x => 351, y => 225),
  (x => 360, y => 225),
  (x => 361, y => 225),
  (x => 362, y => 225),
  (x => 367, y => 225),
  (x => 368, y => 225),
  (x => 369, y => 225),
  (x => 370, y => 225),
  (x => 209, y => 226),
  (x => 210, y => 226),
  (x => 211, y => 226),
  (x => 212, y => 226),
  (x => 213, y => 226),
  (x => 214, y => 226),
  (x => 215, y => 226),
  (x => 216, y => 226),
  (x => 217, y => 226),
  (x => 218, y => 226),
  (x => 219, y => 226),
  (x => 220, y => 226),
  (x => 221, y => 226),
  (x => 222, y => 226),
  (x => 228, y => 226),
  (x => 229, y => 226),
  (x => 230, y => 226),
  (x => 231, y => 226),
  (x => 312, y => 226),
  (x => 313, y => 226),
  (x => 314, y => 226),
  (x => 315, y => 226),
  (x => 316, y => 226),
  (x => 317, y => 226),
  (x => 335, y => 226),
  (x => 336, y => 226),
  (x => 337, y => 226),
  (x => 347, y => 226),
  (x => 348, y => 226),
  (x => 349, y => 226),
  (x => 350, y => 226),
  (x => 351, y => 226),
  (x => 359, y => 226),
  (x => 360, y => 226),
  (x => 361, y => 226),
  (x => 362, y => 226),
  (x => 368, y => 226),
  (x => 369, y => 226),
  (x => 209, y => 227),
  (x => 210, y => 227),
  (x => 211, y => 227),
  (x => 212, y => 227),
  (x => 217, y => 227),
  (x => 218, y => 227),
  (x => 219, y => 227),
  (x => 220, y => 227),
  (x => 221, y => 227),
  (x => 222, y => 227),
  (x => 228, y => 227),
  (x => 229, y => 227),
  (x => 230, y => 227),
  (x => 231, y => 227),
  (x => 310, y => 227),
  (x => 311, y => 227),
  (x => 312, y => 227),
  (x => 313, y => 227),
  (x => 314, y => 227),
  (x => 315, y => 227),
  (x => 316, y => 227),
  (x => 317, y => 227),
  (x => 335, y => 227),
  (x => 336, y => 227),
  (x => 337, y => 227),
  (x => 338, y => 227),
  (x => 346, y => 227),
  (x => 347, y => 227),
  (x => 348, y => 227),
  (x => 349, y => 227),
  (x => 350, y => 227),
  (x => 351, y => 227),
  (x => 359, y => 227),
  (x => 360, y => 227),
  (x => 361, y => 227),
  (x => 362, y => 227),
  (x => 209, y => 228),
  (x => 210, y => 228),
  (x => 211, y => 228),
  (x => 212, y => 228),
  (x => 219, y => 228),
  (x => 220, y => 228),
  (x => 221, y => 228),
  (x => 222, y => 228),
  (x => 223, y => 228),
  (x => 228, y => 228),
  (x => 229, y => 228),
  (x => 230, y => 228),
  (x => 231, y => 228),
  (x => 310, y => 228),
  (x => 311, y => 228),
  (x => 312, y => 228),
  (x => 313, y => 228),
  (x => 314, y => 228),
  (x => 315, y => 228),
  (x => 316, y => 228),
  (x => 317, y => 228),
  (x => 335, y => 228),
  (x => 336, y => 228),
  (x => 337, y => 228),
  (x => 338, y => 228),
  (x => 346, y => 228),
  (x => 347, y => 228),
  (x => 348, y => 228),
  (x => 349, y => 228),
  (x => 350, y => 228),
  (x => 351, y => 228),
  (x => 359, y => 228),
  (x => 360, y => 228),
  (x => 361, y => 228),
  (x => 209, y => 229),
  (x => 210, y => 229),
  (x => 211, y => 229),
  (x => 212, y => 229),
  (x => 220, y => 229),
  (x => 221, y => 229),
  (x => 222, y => 229),
  (x => 223, y => 229),
  (x => 228, y => 229),
  (x => 229, y => 229),
  (x => 230, y => 229),
  (x => 231, y => 229),
  (x => 310, y => 229),
  (x => 311, y => 229),
  (x => 312, y => 229),
  (x => 315, y => 229),
  (x => 316, y => 229),
  (x => 317, y => 229),
  (x => 335, y => 229),
  (x => 336, y => 229),
  (x => 337, y => 229),
  (x => 338, y => 229),
  (x => 346, y => 229),
  (x => 347, y => 229),
  (x => 348, y => 229),
  (x => 349, y => 229),
  (x => 350, y => 229),
  (x => 351, y => 229),
  (x => 359, y => 229),
  (x => 360, y => 229),
  (x => 361, y => 229),
  (x => 209, y => 230),
  (x => 210, y => 230),
  (x => 211, y => 230),
  (x => 212, y => 230),
  (x => 220, y => 230),
  (x => 221, y => 230),
  (x => 222, y => 230),
  (x => 223, y => 230),
  (x => 228, y => 230),
  (x => 229, y => 230),
  (x => 230, y => 230),
  (x => 231, y => 230),
  (x => 310, y => 230),
  (x => 311, y => 230),
  (x => 315, y => 230),
  (x => 316, y => 230),
  (x => 317, y => 230),
  (x => 335, y => 230),
  (x => 336, y => 230),
  (x => 337, y => 230),
  (x => 338, y => 230),
  (x => 346, y => 230),
  (x => 347, y => 230),
  (x => 350, y => 230),
  (x => 351, y => 230),
  (x => 352, y => 230),
  (x => 359, y => 230),
  (x => 360, y => 230),
  (x => 361, y => 230),
  (x => 209, y => 231),
  (x => 210, y => 231),
  (x => 211, y => 231),
  (x => 212, y => 231),
  (x => 220, y => 231),
  (x => 221, y => 231),
  (x => 222, y => 231),
  (x => 223, y => 231),
  (x => 228, y => 231),
  (x => 229, y => 231),
  (x => 230, y => 231),
  (x => 231, y => 231),
  (x => 242, y => 231),
  (x => 243, y => 231),
  (x => 276, y => 231),
  (x => 277, y => 231),
  (x => 296, y => 231),
  (x => 315, y => 231),
  (x => 316, y => 231),
  (x => 317, y => 231),
  (x => 336, y => 231),
  (x => 337, y => 231),
  (x => 338, y => 231),
  (x => 346, y => 231),
  (x => 347, y => 231),
  (x => 350, y => 231),
  (x => 351, y => 231),
  (x => 352, y => 231),
  (x => 359, y => 231),
  (x => 360, y => 231),
  (x => 361, y => 231),
  (x => 385, y => 231),
  (x => 386, y => 231),
  (x => 399, y => 231),
  (x => 400, y => 231),
  (x => 401, y => 231),
  (x => 209, y => 232),
  (x => 210, y => 232),
  (x => 211, y => 232),
  (x => 212, y => 232),
  (x => 220, y => 232),
  (x => 221, y => 232),
  (x => 222, y => 232),
  (x => 223, y => 232),
  (x => 228, y => 232),
  (x => 229, y => 232),
  (x => 230, y => 232),
  (x => 231, y => 232),
  (x => 238, y => 232),
  (x => 239, y => 232),
  (x => 240, y => 232),
  (x => 241, y => 232),
  (x => 242, y => 232),
  (x => 243, y => 232),
  (x => 244, y => 232),
  (x => 245, y => 232),
  (x => 246, y => 232),
  (x => 252, y => 232),
  (x => 253, y => 232),
  (x => 254, y => 232),
  (x => 255, y => 232),
  (x => 264, y => 232),
  (x => 265, y => 232),
  (x => 266, y => 232),
  (x => 267, y => 232),
  (x => 274, y => 232),
  (x => 275, y => 232),
  (x => 276, y => 232),
  (x => 277, y => 232),
  (x => 278, y => 232),
  (x => 279, y => 232),
  (x => 280, y => 232),
  (x => 288, y => 232),
  (x => 289, y => 232),
  (x => 290, y => 232),
  (x => 291, y => 232),
  (x => 294, y => 232),
  (x => 295, y => 232),
  (x => 296, y => 232),
  (x => 315, y => 232),
  (x => 316, y => 232),
  (x => 317, y => 232),
  (x => 336, y => 232),
  (x => 337, y => 232),
  (x => 338, y => 232),
  (x => 345, y => 232),
  (x => 346, y => 232),
  (x => 347, y => 232),
  (x => 350, y => 232),
  (x => 351, y => 232),
  (x => 352, y => 232),
  (x => 358, y => 232),
  (x => 359, y => 232),
  (x => 360, y => 232),
  (x => 361, y => 232),
  (x => 367, y => 232),
  (x => 368, y => 232),
  (x => 369, y => 232),
  (x => 370, y => 232),
  (x => 376, y => 232),
  (x => 377, y => 232),
  (x => 378, y => 232),
  (x => 379, y => 232),
  (x => 383, y => 232),
  (x => 384, y => 232),
  (x => 385, y => 232),
  (x => 386, y => 232),
  (x => 387, y => 232),
  (x => 397, y => 232),
  (x => 398, y => 232),
  (x => 399, y => 232),
  (x => 400, y => 232),
  (x => 401, y => 232),
  (x => 402, y => 232),
  (x => 403, y => 232),
  (x => 209, y => 233),
  (x => 210, y => 233),
  (x => 211, y => 233),
  (x => 212, y => 233),
  (x => 220, y => 233),
  (x => 221, y => 233),
  (x => 222, y => 233),
  (x => 223, y => 233),
  (x => 228, y => 233),
  (x => 229, y => 233),
  (x => 230, y => 233),
  (x => 231, y => 233),
  (x => 238, y => 233),
  (x => 239, y => 233),
  (x => 240, y => 233),
  (x => 241, y => 233),
  (x => 242, y => 233),
  (x => 243, y => 233),
  (x => 244, y => 233),
  (x => 245, y => 233),
  (x => 246, y => 233),
  (x => 247, y => 233),
  (x => 253, y => 233),
  (x => 254, y => 233),
  (x => 255, y => 233),
  (x => 256, y => 233),
  (x => 264, y => 233),
  (x => 265, y => 233),
  (x => 266, y => 233),
  (x => 273, y => 233),
  (x => 274, y => 233),
  (x => 275, y => 233),
  (x => 276, y => 233),
  (x => 277, y => 233),
  (x => 278, y => 233),
  (x => 279, y => 233),
  (x => 280, y => 233),
  (x => 281, y => 233),
  (x => 288, y => 233),
  (x => 289, y => 233),
  (x => 290, y => 233),
  (x => 294, y => 233),
  (x => 295, y => 233),
  (x => 296, y => 233),
  (x => 315, y => 233),
  (x => 316, y => 233),
  (x => 317, y => 233),
  (x => 336, y => 233),
  (x => 337, y => 233),
  (x => 338, y => 233),
  (x => 339, y => 233),
  (x => 345, y => 233),
  (x => 346, y => 233),
  (x => 347, y => 233),
  (x => 350, y => 233),
  (x => 351, y => 233),
  (x => 352, y => 233),
  (x => 358, y => 233),
  (x => 359, y => 233),
  (x => 360, y => 233),
  (x => 367, y => 233),
  (x => 368, y => 233),
  (x => 369, y => 233),
  (x => 370, y => 233),
  (x => 376, y => 233),
  (x => 377, y => 233),
  (x => 378, y => 233),
  (x => 379, y => 233),
  (x => 382, y => 233),
  (x => 383, y => 233),
  (x => 384, y => 233),
  (x => 385, y => 233),
  (x => 386, y => 233),
  (x => 387, y => 233),
  (x => 388, y => 233),
  (x => 396, y => 233),
  (x => 397, y => 233),
  (x => 398, y => 233),
  (x => 399, y => 233),
  (x => 400, y => 233),
  (x => 401, y => 233),
  (x => 402, y => 233),
  (x => 403, y => 233),
  (x => 209, y => 234),
  (x => 210, y => 234),
  (x => 211, y => 234),
  (x => 212, y => 234),
  (x => 220, y => 234),
  (x => 221, y => 234),
  (x => 222, y => 234),
  (x => 223, y => 234),
  (x => 228, y => 234),
  (x => 229, y => 234),
  (x => 230, y => 234),
  (x => 231, y => 234),
  (x => 238, y => 234),
  (x => 239, y => 234),
  (x => 240, y => 234),
  (x => 241, y => 234),
  (x => 243, y => 234),
  (x => 244, y => 234),
  (x => 245, y => 234),
  (x => 246, y => 234),
  (x => 247, y => 234),
  (x => 253, y => 234),
  (x => 254, y => 234),
  (x => 255, y => 234),
  (x => 256, y => 234),
  (x => 264, y => 234),
  (x => 265, y => 234),
  (x => 266, y => 234),
  (x => 272, y => 234),
  (x => 273, y => 234),
  (x => 274, y => 234),
  (x => 275, y => 234),
  (x => 276, y => 234),
  (x => 278, y => 234),
  (x => 279, y => 234),
  (x => 280, y => 234),
  (x => 281, y => 234),
  (x => 288, y => 234),
  (x => 289, y => 234),
  (x => 290, y => 234),
  (x => 293, y => 234),
  (x => 294, y => 234),
  (x => 295, y => 234),
  (x => 296, y => 234),
  (x => 315, y => 234),
  (x => 316, y => 234),
  (x => 317, y => 234),
  (x => 336, y => 234),
  (x => 337, y => 234),
  (x => 338, y => 234),
  (x => 339, y => 234),
  (x => 345, y => 234),
  (x => 346, y => 234),
  (x => 350, y => 234),
  (x => 351, y => 234),
  (x => 352, y => 234),
  (x => 358, y => 234),
  (x => 359, y => 234),
  (x => 360, y => 234),
  (x => 367, y => 234),
  (x => 368, y => 234),
  (x => 369, y => 234),
  (x => 370, y => 234),
  (x => 376, y => 234),
  (x => 377, y => 234),
  (x => 378, y => 234),
  (x => 379, y => 234),
  (x => 382, y => 234),
  (x => 383, y => 234),
  (x => 384, y => 234),
  (x => 385, y => 234),
  (x => 386, y => 234),
  (x => 387, y => 234),
  (x => 388, y => 234),
  (x => 389, y => 234),
  (x => 395, y => 234),
  (x => 396, y => 234),
  (x => 397, y => 234),
  (x => 398, y => 234),
  (x => 399, y => 234),
  (x => 400, y => 234),
  (x => 401, y => 234),
  (x => 402, y => 234),
  (x => 403, y => 234),
  (x => 209, y => 235),
  (x => 210, y => 235),
  (x => 211, y => 235),
  (x => 212, y => 235),
  (x => 220, y => 235),
  (x => 221, y => 235),
  (x => 222, y => 235),
  (x => 223, y => 235),
  (x => 228, y => 235),
  (x => 229, y => 235),
  (x => 230, y => 235),
  (x => 231, y => 235),
  (x => 238, y => 235),
  (x => 245, y => 235),
  (x => 246, y => 235),
  (x => 247, y => 235),
  (x => 254, y => 235),
  (x => 255, y => 235),
  (x => 256, y => 235),
  (x => 264, y => 235),
  (x => 265, y => 235),
  (x => 266, y => 235),
  (x => 272, y => 235),
  (x => 273, y => 235),
  (x => 274, y => 235),
  (x => 280, y => 235),
  (x => 281, y => 235),
  (x => 282, y => 235),
  (x => 288, y => 235),
  (x => 289, y => 235),
  (x => 290, y => 235),
  (x => 291, y => 235),
  (x => 292, y => 235),
  (x => 293, y => 235),
  (x => 294, y => 235),
  (x => 295, y => 235),
  (x => 296, y => 235),
  (x => 315, y => 235),
  (x => 316, y => 235),
  (x => 317, y => 235),
  (x => 337, y => 235),
  (x => 338, y => 235),
  (x => 339, y => 235),
  (x => 345, y => 235),
  (x => 346, y => 235),
  (x => 350, y => 235),
  (x => 351, y => 235),
  (x => 352, y => 235),
  (x => 358, y => 235),
  (x => 359, y => 235),
  (x => 360, y => 235),
  (x => 367, y => 235),
  (x => 368, y => 235),
  (x => 369, y => 235),
  (x => 370, y => 235),
  (x => 376, y => 235),
  (x => 377, y => 235),
  (x => 378, y => 235),
  (x => 379, y => 235),
  (x => 380, y => 235),
  (x => 381, y => 235),
  (x => 385, y => 235),
  (x => 386, y => 235),
  (x => 387, y => 235),
  (x => 388, y => 235),
  (x => 389, y => 235),
  (x => 395, y => 235),
  (x => 396, y => 235),
  (x => 397, y => 235),
  (x => 209, y => 236),
  (x => 210, y => 236),
  (x => 211, y => 236),
  (x => 212, y => 236),
  (x => 219, y => 236),
  (x => 220, y => 236),
  (x => 221, y => 236),
  (x => 222, y => 236),
  (x => 228, y => 236),
  (x => 229, y => 236),
  (x => 230, y => 236),
  (x => 231, y => 236),
  (x => 246, y => 236),
  (x => 247, y => 236),
  (x => 248, y => 236),
  (x => 254, y => 236),
  (x => 255, y => 236),
  (x => 256, y => 236),
  (x => 263, y => 236),
  (x => 264, y => 236),
  (x => 265, y => 236),
  (x => 271, y => 236),
  (x => 272, y => 236),
  (x => 273, y => 236),
  (x => 280, y => 236),
  (x => 281, y => 236),
  (x => 282, y => 236),
  (x => 288, y => 236),
  (x => 289, y => 236),
  (x => 290, y => 236),
  (x => 291, y => 236),
  (x => 292, y => 236),
  (x => 315, y => 236),
  (x => 316, y => 236),
  (x => 317, y => 236),
  (x => 337, y => 236),
  (x => 338, y => 236),
  (x => 339, y => 236),
  (x => 345, y => 236),
  (x => 346, y => 236),
  (x => 351, y => 236),
  (x => 352, y => 236),
  (x => 353, y => 236),
  (x => 358, y => 236),
  (x => 359, y => 236),
  (x => 360, y => 236),
  (x => 367, y => 236),
  (x => 368, y => 236),
  (x => 369, y => 236),
  (x => 370, y => 236),
  (x => 376, y => 236),
  (x => 377, y => 236),
  (x => 378, y => 236),
  (x => 379, y => 236),
  (x => 380, y => 236),
  (x => 386, y => 236),
  (x => 387, y => 236),
  (x => 388, y => 236),
  (x => 389, y => 236),
  (x => 394, y => 236),
  (x => 395, y => 236),
  (x => 396, y => 236),
  (x => 397, y => 236),
  (x => 209, y => 237),
  (x => 210, y => 237),
  (x => 211, y => 237),
  (x => 212, y => 237),
  (x => 218, y => 237),
  (x => 219, y => 237),
  (x => 220, y => 237),
  (x => 221, y => 237),
  (x => 222, y => 237),
  (x => 228, y => 237),
  (x => 229, y => 237),
  (x => 230, y => 237),
  (x => 231, y => 237),
  (x => 246, y => 237),
  (x => 247, y => 237),
  (x => 248, y => 237),
  (x => 254, y => 237),
  (x => 255, y => 237),
  (x => 256, y => 237),
  (x => 263, y => 237),
  (x => 264, y => 237),
  (x => 265, y => 237),
  (x => 271, y => 237),
  (x => 272, y => 237),
  (x => 273, y => 237),
  (x => 281, y => 237),
  (x => 282, y => 237),
  (x => 288, y => 237),
  (x => 289, y => 237),
  (x => 290, y => 237),
  (x => 291, y => 237),
  (x => 315, y => 237),
  (x => 316, y => 237),
  (x => 317, y => 237),
  (x => 337, y => 237),
  (x => 338, y => 237),
  (x => 339, y => 237),
  (x => 344, y => 237),
  (x => 345, y => 237),
  (x => 346, y => 237),
  (x => 351, y => 237),
  (x => 352, y => 237),
  (x => 353, y => 237),
  (x => 358, y => 237),
  (x => 359, y => 237),
  (x => 360, y => 237),
  (x => 367, y => 237),
  (x => 368, y => 237),
  (x => 369, y => 237),
  (x => 370, y => 237),
  (x => 376, y => 237),
  (x => 377, y => 237),
  (x => 378, y => 237),
  (x => 379, y => 237),
  (x => 386, y => 237),
  (x => 387, y => 237),
  (x => 388, y => 237),
  (x => 389, y => 237),
  (x => 394, y => 237),
  (x => 395, y => 237),
  (x => 396, y => 237),
  (x => 397, y => 237),
  (x => 209, y => 238),
  (x => 210, y => 238),
  (x => 211, y => 238),
  (x => 212, y => 238),
  (x => 213, y => 238),
  (x => 214, y => 238),
  (x => 215, y => 238),
  (x => 216, y => 238),
  (x => 217, y => 238),
  (x => 218, y => 238),
  (x => 219, y => 238),
  (x => 220, y => 238),
  (x => 221, y => 238),
  (x => 228, y => 238),
  (x => 229, y => 238),
  (x => 230, y => 238),
  (x => 231, y => 238),
  (x => 246, y => 238),
  (x => 247, y => 238),
  (x => 248, y => 238),
  (x => 254, y => 238),
  (x => 255, y => 238),
  (x => 256, y => 238),
  (x => 257, y => 238),
  (x => 263, y => 238),
  (x => 264, y => 238),
  (x => 265, y => 238),
  (x => 271, y => 238),
  (x => 272, y => 238),
  (x => 273, y => 238),
  (x => 281, y => 238),
  (x => 282, y => 238),
  (x => 283, y => 238),
  (x => 288, y => 238),
  (x => 289, y => 238),
  (x => 290, y => 238),
  (x => 291, y => 238),
  (x => 315, y => 238),
  (x => 316, y => 238),
  (x => 317, y => 238),
  (x => 337, y => 238),
  (x => 338, y => 238),
  (x => 339, y => 238),
  (x => 344, y => 238),
  (x => 345, y => 238),
  (x => 346, y => 238),
  (x => 351, y => 238),
  (x => 352, y => 238),
  (x => 353, y => 238),
  (x => 358, y => 238),
  (x => 359, y => 238),
  (x => 367, y => 238),
  (x => 368, y => 238),
  (x => 369, y => 238),
  (x => 370, y => 238),
  (x => 376, y => 238),
  (x => 377, y => 238),
  (x => 378, y => 238),
  (x => 379, y => 238),
  (x => 387, y => 238),
  (x => 388, y => 238),
  (x => 389, y => 238),
  (x => 394, y => 238),
  (x => 395, y => 238),
  (x => 396, y => 238),
  (x => 397, y => 238),
  (x => 209, y => 239),
  (x => 210, y => 239),
  (x => 211, y => 239),
  (x => 212, y => 239),
  (x => 213, y => 239),
  (x => 214, y => 239),
  (x => 215, y => 239),
  (x => 216, y => 239),
  (x => 217, y => 239),
  (x => 218, y => 239),
  (x => 219, y => 239),
  (x => 220, y => 239),
  (x => 221, y => 239),
  (x => 228, y => 239),
  (x => 229, y => 239),
  (x => 230, y => 239),
  (x => 231, y => 239),
  (x => 244, y => 239),
  (x => 245, y => 239),
  (x => 246, y => 239),
  (x => 247, y => 239),
  (x => 248, y => 239),
  (x => 255, y => 239),
  (x => 256, y => 239),
  (x => 257, y => 239),
  (x => 263, y => 239),
  (x => 264, y => 239),
  (x => 270, y => 239),
  (x => 271, y => 239),
  (x => 272, y => 239),
  (x => 273, y => 239),
  (x => 281, y => 239),
  (x => 282, y => 239),
  (x => 283, y => 239),
  (x => 288, y => 239),
  (x => 289, y => 239),
  (x => 290, y => 239),
  (x => 291, y => 239),
  (x => 315, y => 239),
  (x => 316, y => 239),
  (x => 317, y => 239),
  (x => 337, y => 239),
  (x => 338, y => 239),
  (x => 339, y => 239),
  (x => 340, y => 239),
  (x => 344, y => 239),
  (x => 345, y => 239),
  (x => 346, y => 239),
  (x => 351, y => 239),
  (x => 352, y => 239),
  (x => 353, y => 239),
  (x => 357, y => 239),
  (x => 358, y => 239),
  (x => 359, y => 239),
  (x => 367, y => 239),
  (x => 368, y => 239),
  (x => 369, y => 239),
  (x => 370, y => 239),
  (x => 376, y => 239),
  (x => 377, y => 239),
  (x => 378, y => 239),
  (x => 379, y => 239),
  (x => 387, y => 239),
  (x => 388, y => 239),
  (x => 389, y => 239),
  (x => 395, y => 239),
  (x => 396, y => 239),
  (x => 397, y => 239),
  (x => 398, y => 239),
  (x => 399, y => 239),
  (x => 209, y => 240),
  (x => 210, y => 240),
  (x => 211, y => 240),
  (x => 212, y => 240),
  (x => 213, y => 240),
  (x => 214, y => 240),
  (x => 215, y => 240),
  (x => 216, y => 240),
  (x => 217, y => 240),
  (x => 218, y => 240),
  (x => 219, y => 240),
  (x => 228, y => 240),
  (x => 229, y => 240),
  (x => 230, y => 240),
  (x => 231, y => 240),
  (x => 239, y => 240),
  (x => 240, y => 240),
  (x => 241, y => 240),
  (x => 242, y => 240),
  (x => 243, y => 240),
  (x => 244, y => 240),
  (x => 245, y => 240),
  (x => 246, y => 240),
  (x => 247, y => 240),
  (x => 248, y => 240),
  (x => 255, y => 240),
  (x => 256, y => 240),
  (x => 257, y => 240),
  (x => 262, y => 240),
  (x => 263, y => 240),
  (x => 264, y => 240),
  (x => 270, y => 240),
  (x => 271, y => 240),
  (x => 272, y => 240),
  (x => 273, y => 240),
  (x => 274, y => 240),
  (x => 275, y => 240),
  (x => 276, y => 240),
  (x => 277, y => 240),
  (x => 278, y => 240),
  (x => 279, y => 240),
  (x => 280, y => 240),
  (x => 281, y => 240),
  (x => 282, y => 240),
  (x => 283, y => 240),
  (x => 288, y => 240),
  (x => 289, y => 240),
  (x => 290, y => 240),
  (x => 315, y => 240),
  (x => 316, y => 240),
  (x => 317, y => 240),
  (x => 338, y => 240),
  (x => 339, y => 240),
  (x => 340, y => 240),
  (x => 344, y => 240),
  (x => 345, y => 240),
  (x => 351, y => 240),
  (x => 352, y => 240),
  (x => 353, y => 240),
  (x => 357, y => 240),
  (x => 358, y => 240),
  (x => 359, y => 240),
  (x => 367, y => 240),
  (x => 368, y => 240),
  (x => 369, y => 240),
  (x => 370, y => 240),
  (x => 376, y => 240),
  (x => 377, y => 240),
  (x => 378, y => 240),
  (x => 379, y => 240),
  (x => 387, y => 240),
  (x => 388, y => 240),
  (x => 389, y => 240),
  (x => 395, y => 240),
  (x => 396, y => 240),
  (x => 397, y => 240),
  (x => 398, y => 240),
  (x => 399, y => 240),
  (x => 400, y => 240),
  (x => 401, y => 240),
  (x => 209, y => 241),
  (x => 210, y => 241),
  (x => 211, y => 241),
  (x => 212, y => 241),
  (x => 213, y => 241),
  (x => 214, y => 241),
  (x => 215, y => 241),
  (x => 216, y => 241),
  (x => 217, y => 241),
  (x => 228, y => 241),
  (x => 229, y => 241),
  (x => 230, y => 241),
  (x => 231, y => 241),
  (x => 238, y => 241),
  (x => 239, y => 241),
  (x => 240, y => 241),
  (x => 241, y => 241),
  (x => 242, y => 241),
  (x => 243, y => 241),
  (x => 244, y => 241),
  (x => 245, y => 241),
  (x => 246, y => 241),
  (x => 247, y => 241),
  (x => 248, y => 241),
  (x => 255, y => 241),
  (x => 256, y => 241),
  (x => 257, y => 241),
  (x => 262, y => 241),
  (x => 263, y => 241),
  (x => 264, y => 241),
  (x => 270, y => 241),
  (x => 271, y => 241),
  (x => 272, y => 241),
  (x => 273, y => 241),
  (x => 274, y => 241),
  (x => 275, y => 241),
  (x => 276, y => 241),
  (x => 277, y => 241),
  (x => 278, y => 241),
  (x => 279, y => 241),
  (x => 280, y => 241),
  (x => 281, y => 241),
  (x => 282, y => 241),
  (x => 283, y => 241),
  (x => 288, y => 241),
  (x => 289, y => 241),
  (x => 290, y => 241),
  (x => 315, y => 241),
  (x => 316, y => 241),
  (x => 317, y => 241),
  (x => 338, y => 241),
  (x => 339, y => 241),
  (x => 340, y => 241),
  (x => 344, y => 241),
  (x => 345, y => 241),
  (x => 352, y => 241),
  (x => 353, y => 241),
  (x => 354, y => 241),
  (x => 357, y => 241),
  (x => 358, y => 241),
  (x => 359, y => 241),
  (x => 367, y => 241),
  (x => 368, y => 241),
  (x => 369, y => 241),
  (x => 370, y => 241),
  (x => 376, y => 241),
  (x => 377, y => 241),
  (x => 378, y => 241),
  (x => 379, y => 241),
  (x => 387, y => 241),
  (x => 388, y => 241),
  (x => 389, y => 241),
  (x => 396, y => 241),
  (x => 397, y => 241),
  (x => 398, y => 241),
  (x => 399, y => 241),
  (x => 400, y => 241),
  (x => 401, y => 241),
  (x => 402, y => 241),
  (x => 209, y => 242),
  (x => 210, y => 242),
  (x => 211, y => 242),
  (x => 212, y => 242),
  (x => 228, y => 242),
  (x => 229, y => 242),
  (x => 230, y => 242),
  (x => 231, y => 242),
  (x => 237, y => 242),
  (x => 238, y => 242),
  (x => 239, y => 242),
  (x => 240, y => 242),
  (x => 246, y => 242),
  (x => 247, y => 242),
  (x => 248, y => 242),
  (x => 256, y => 242),
  (x => 257, y => 242),
  (x => 258, y => 242),
  (x => 262, y => 242),
  (x => 263, y => 242),
  (x => 264, y => 242),
  (x => 270, y => 242),
  (x => 271, y => 242),
  (x => 272, y => 242),
  (x => 273, y => 242),
  (x => 274, y => 242),
  (x => 275, y => 242),
  (x => 276, y => 242),
  (x => 277, y => 242),
  (x => 278, y => 242),
  (x => 279, y => 242),
  (x => 280, y => 242),
  (x => 281, y => 242),
  (x => 282, y => 242),
  (x => 283, y => 242),
  (x => 288, y => 242),
  (x => 289, y => 242),
  (x => 290, y => 242),
  (x => 315, y => 242),
  (x => 316, y => 242),
  (x => 317, y => 242),
  (x => 338, y => 242),
  (x => 339, y => 242),
  (x => 340, y => 242),
  (x => 343, y => 242),
  (x => 344, y => 242),
  (x => 345, y => 242),
  (x => 352, y => 242),
  (x => 353, y => 242),
  (x => 354, y => 242),
  (x => 357, y => 242),
  (x => 358, y => 242),
  (x => 359, y => 242),
  (x => 367, y => 242),
  (x => 368, y => 242),
  (x => 369, y => 242),
  (x => 370, y => 242),
  (x => 376, y => 242),
  (x => 377, y => 242),
  (x => 378, y => 242),
  (x => 379, y => 242),
  (x => 387, y => 242),
  (x => 388, y => 242),
  (x => 389, y => 242),
  (x => 397, y => 242),
  (x => 398, y => 242),
  (x => 399, y => 242),
  (x => 400, y => 242),
  (x => 401, y => 242),
  (x => 402, y => 242),
  (x => 403, y => 242),
  (x => 209, y => 243),
  (x => 210, y => 243),
  (x => 211, y => 243),
  (x => 212, y => 243),
  (x => 228, y => 243),
  (x => 229, y => 243),
  (x => 230, y => 243),
  (x => 231, y => 243),
  (x => 237, y => 243),
  (x => 238, y => 243),
  (x => 239, y => 243),
  (x => 246, y => 243),
  (x => 247, y => 243),
  (x => 248, y => 243),
  (x => 256, y => 243),
  (x => 257, y => 243),
  (x => 258, y => 243),
  (x => 262, y => 243),
  (x => 263, y => 243),
  (x => 270, y => 243),
  (x => 271, y => 243),
  (x => 272, y => 243),
  (x => 273, y => 243),
  (x => 288, y => 243),
  (x => 289, y => 243),
  (x => 290, y => 243),
  (x => 315, y => 243),
  (x => 316, y => 243),
  (x => 317, y => 243),
  (x => 338, y => 243),
  (x => 339, y => 243),
  (x => 340, y => 243),
  (x => 343, y => 243),
  (x => 344, y => 243),
  (x => 345, y => 243),
  (x => 352, y => 243),
  (x => 353, y => 243),
  (x => 354, y => 243),
  (x => 357, y => 243),
  (x => 358, y => 243),
  (x => 367, y => 243),
  (x => 368, y => 243),
  (x => 369, y => 243),
  (x => 370, y => 243),
  (x => 376, y => 243),
  (x => 377, y => 243),
  (x => 378, y => 243),
  (x => 379, y => 243),
  (x => 387, y => 243),
  (x => 388, y => 243),
  (x => 389, y => 243),
  (x => 399, y => 243),
  (x => 400, y => 243),
  (x => 401, y => 243),
  (x => 402, y => 243),
  (x => 403, y => 243),
  (x => 404, y => 243),
  (x => 209, y => 244),
  (x => 210, y => 244),
  (x => 211, y => 244),
  (x => 212, y => 244),
  (x => 228, y => 244),
  (x => 229, y => 244),
  (x => 230, y => 244),
  (x => 231, y => 244),
  (x => 236, y => 244),
  (x => 237, y => 244),
  (x => 238, y => 244),
  (x => 246, y => 244),
  (x => 247, y => 244),
  (x => 248, y => 244),
  (x => 256, y => 244),
  (x => 257, y => 244),
  (x => 258, y => 244),
  (x => 261, y => 244),
  (x => 262, y => 244),
  (x => 263, y => 244),
  (x => 270, y => 244),
  (x => 271, y => 244),
  (x => 272, y => 244),
  (x => 273, y => 244),
  (x => 288, y => 244),
  (x => 289, y => 244),
  (x => 290, y => 244),
  (x => 315, y => 244),
  (x => 316, y => 244),
  (x => 317, y => 244),
  (x => 338, y => 244),
  (x => 339, y => 244),
  (x => 340, y => 244),
  (x => 343, y => 244),
  (x => 344, y => 244),
  (x => 345, y => 244),
  (x => 352, y => 244),
  (x => 353, y => 244),
  (x => 354, y => 244),
  (x => 357, y => 244),
  (x => 358, y => 244),
  (x => 367, y => 244),
  (x => 368, y => 244),
  (x => 369, y => 244),
  (x => 370, y => 244),
  (x => 376, y => 244),
  (x => 377, y => 244),
  (x => 378, y => 244),
  (x => 379, y => 244),
  (x => 387, y => 244),
  (x => 388, y => 244),
  (x => 389, y => 244),
  (x => 401, y => 244),
  (x => 402, y => 244),
  (x => 403, y => 244),
  (x => 404, y => 244),
  (x => 209, y => 245),
  (x => 210, y => 245),
  (x => 211, y => 245),
  (x => 212, y => 245),
  (x => 228, y => 245),
  (x => 229, y => 245),
  (x => 230, y => 245),
  (x => 231, y => 245),
  (x => 236, y => 245),
  (x => 237, y => 245),
  (x => 238, y => 245),
  (x => 246, y => 245),
  (x => 247, y => 245),
  (x => 248, y => 245),
  (x => 257, y => 245),
  (x => 258, y => 245),
  (x => 261, y => 245),
  (x => 262, y => 245),
  (x => 263, y => 245),
  (x => 271, y => 245),
  (x => 272, y => 245),
  (x => 273, y => 245),
  (x => 288, y => 245),
  (x => 289, y => 245),
  (x => 290, y => 245),
  (x => 315, y => 245),
  (x => 316, y => 245),
  (x => 317, y => 245),
  (x => 338, y => 245),
  (x => 339, y => 245),
  (x => 340, y => 245),
  (x => 343, y => 245),
  (x => 344, y => 245),
  (x => 352, y => 245),
  (x => 353, y => 245),
  (x => 354, y => 245),
  (x => 357, y => 245),
  (x => 358, y => 245),
  (x => 367, y => 245),
  (x => 368, y => 245),
  (x => 369, y => 245),
  (x => 370, y => 245),
  (x => 376, y => 245),
  (x => 377, y => 245),
  (x => 378, y => 245),
  (x => 379, y => 245),
  (x => 387, y => 245),
  (x => 388, y => 245),
  (x => 389, y => 245),
  (x => 402, y => 245),
  (x => 403, y => 245),
  (x => 404, y => 245),
  (x => 209, y => 246),
  (x => 210, y => 246),
  (x => 211, y => 246),
  (x => 212, y => 246),
  (x => 228, y => 246),
  (x => 229, y => 246),
  (x => 230, y => 246),
  (x => 231, y => 246),
  (x => 236, y => 246),
  (x => 237, y => 246),
  (x => 238, y => 246),
  (x => 245, y => 246),
  (x => 246, y => 246),
  (x => 247, y => 246),
  (x => 248, y => 246),
  (x => 257, y => 246),
  (x => 258, y => 246),
  (x => 261, y => 246),
  (x => 262, y => 246),
  (x => 271, y => 246),
  (x => 272, y => 246),
  (x => 273, y => 246),
  (x => 288, y => 246),
  (x => 289, y => 246),
  (x => 290, y => 246),
  (x => 315, y => 246),
  (x => 316, y => 246),
  (x => 317, y => 246),
  (x => 339, y => 246),
  (x => 340, y => 246),
  (x => 341, y => 246),
  (x => 342, y => 246),
  (x => 343, y => 246),
  (x => 344, y => 246),
  (x => 353, y => 246),
  (x => 354, y => 246),
  (x => 355, y => 246),
  (x => 356, y => 246),
  (x => 357, y => 246),
  (x => 358, y => 246),
  (x => 367, y => 246),
  (x => 368, y => 246),
  (x => 369, y => 246),
  (x => 370, y => 246),
  (x => 376, y => 246),
  (x => 377, y => 246),
  (x => 378, y => 246),
  (x => 379, y => 246),
  (x => 387, y => 246),
  (x => 388, y => 246),
  (x => 389, y => 246),
  (x => 402, y => 246),
  (x => 403, y => 246),
  (x => 404, y => 246),
  (x => 209, y => 247),
  (x => 210, y => 247),
  (x => 211, y => 247),
  (x => 212, y => 247),
  (x => 228, y => 247),
  (x => 229, y => 247),
  (x => 230, y => 247),
  (x => 231, y => 247),
  (x => 236, y => 247),
  (x => 237, y => 247),
  (x => 238, y => 247),
  (x => 239, y => 247),
  (x => 245, y => 247),
  (x => 246, y => 247),
  (x => 247, y => 247),
  (x => 248, y => 247),
  (x => 257, y => 247),
  (x => 258, y => 247),
  (x => 259, y => 247),
  (x => 260, y => 247),
  (x => 261, y => 247),
  (x => 262, y => 247),
  (x => 271, y => 247),
  (x => 272, y => 247),
  (x => 273, y => 247),
  (x => 274, y => 247),
  (x => 288, y => 247),
  (x => 289, y => 247),
  (x => 290, y => 247),
  (x => 315, y => 247),
  (x => 316, y => 247),
  (x => 317, y => 247),
  (x => 339, y => 247),
  (x => 340, y => 247),
  (x => 341, y => 247),
  (x => 342, y => 247),
  (x => 343, y => 247),
  (x => 344, y => 247),
  (x => 353, y => 247),
  (x => 354, y => 247),
  (x => 355, y => 247),
  (x => 356, y => 247),
  (x => 357, y => 247),
  (x => 358, y => 247),
  (x => 367, y => 247),
  (x => 368, y => 247),
  (x => 369, y => 247),
  (x => 370, y => 247),
  (x => 376, y => 247),
  (x => 377, y => 247),
  (x => 378, y => 247),
  (x => 379, y => 247),
  (x => 387, y => 247),
  (x => 388, y => 247),
  (x => 389, y => 247),
  (x => 402, y => 247),
  (x => 403, y => 247),
  (x => 404, y => 247),
  (x => 209, y => 248),
  (x => 210, y => 248),
  (x => 211, y => 248),
  (x => 212, y => 248),
  (x => 228, y => 248),
  (x => 229, y => 248),
  (x => 230, y => 248),
  (x => 231, y => 248),
  (x => 236, y => 248),
  (x => 237, y => 248),
  (x => 238, y => 248),
  (x => 239, y => 248),
  (x => 240, y => 248),
  (x => 243, y => 248),
  (x => 244, y => 248),
  (x => 245, y => 248),
  (x => 246, y => 248),
  (x => 247, y => 248),
  (x => 248, y => 248),
  (x => 257, y => 248),
  (x => 258, y => 248),
  (x => 259, y => 248),
  (x => 260, y => 248),
  (x => 261, y => 248),
  (x => 262, y => 248),
  (x => 272, y => 248),
  (x => 273, y => 248),
  (x => 274, y => 248),
  (x => 275, y => 248),
  (x => 276, y => 248),
  (x => 281, y => 248),
  (x => 288, y => 248),
  (x => 289, y => 248),
  (x => 290, y => 248),
  (x => 315, y => 248),
  (x => 316, y => 248),
  (x => 317, y => 248),
  (x => 339, y => 248),
  (x => 340, y => 248),
  (x => 341, y => 248),
  (x => 342, y => 248),
  (x => 343, y => 248),
  (x => 344, y => 248),
  (x => 353, y => 248),
  (x => 354, y => 248),
  (x => 355, y => 248),
  (x => 356, y => 248),
  (x => 357, y => 248),
  (x => 367, y => 248),
  (x => 368, y => 248),
  (x => 369, y => 248),
  (x => 370, y => 248),
  (x => 376, y => 248),
  (x => 377, y => 248),
  (x => 378, y => 248),
  (x => 379, y => 248),
  (x => 387, y => 248),
  (x => 388, y => 248),
  (x => 389, y => 248),
  (x => 394, y => 248),
  (x => 395, y => 248),
  (x => 401, y => 248),
  (x => 402, y => 248),
  (x => 403, y => 248),
  (x => 404, y => 248),
  (x => 209, y => 249),
  (x => 210, y => 249),
  (x => 211, y => 249),
  (x => 212, y => 249),
  (x => 228, y => 249),
  (x => 229, y => 249),
  (x => 230, y => 249),
  (x => 231, y => 249),
  (x => 237, y => 249),
  (x => 238, y => 249),
  (x => 239, y => 249),
  (x => 240, y => 249),
  (x => 241, y => 249),
  (x => 242, y => 249),
  (x => 243, y => 249),
  (x => 246, y => 249),
  (x => 247, y => 249),
  (x => 248, y => 249),
  (x => 258, y => 249),
  (x => 259, y => 249),
  (x => 260, y => 249),
  (x => 261, y => 249),
  (x => 262, y => 249),
  (x => 272, y => 249),
  (x => 273, y => 249),
  (x => 274, y => 249),
  (x => 275, y => 249),
  (x => 276, y => 249),
  (x => 277, y => 249),
  (x => 278, y => 249),
  (x => 279, y => 249),
  (x => 280, y => 249),
  (x => 281, y => 249),
  (x => 288, y => 249),
  (x => 289, y => 249),
  (x => 290, y => 249),
  (x => 315, y => 249),
  (x => 316, y => 249),
  (x => 317, y => 249),
  (x => 339, y => 249),
  (x => 340, y => 249),
  (x => 341, y => 249),
  (x => 342, y => 249),
  (x => 343, y => 249),
  (x => 353, y => 249),
  (x => 354, y => 249),
  (x => 355, y => 249),
  (x => 356, y => 249),
  (x => 357, y => 249),
  (x => 367, y => 249),
  (x => 368, y => 249),
  (x => 369, y => 249),
  (x => 370, y => 249),
  (x => 376, y => 249),
  (x => 377, y => 249),
  (x => 378, y => 249),
  (x => 379, y => 249),
  (x => 387, y => 249),
  (x => 388, y => 249),
  (x => 389, y => 249),
  (x => 394, y => 249),
  (x => 395, y => 249),
  (x => 396, y => 249),
  (x => 397, y => 249),
  (x => 398, y => 249),
  (x => 399, y => 249),
  (x => 400, y => 249),
  (x => 401, y => 249),
  (x => 402, y => 249),
  (x => 403, y => 249),
  (x => 209, y => 250),
  (x => 210, y => 250),
  (x => 211, y => 250),
  (x => 212, y => 250),
  (x => 228, y => 250),
  (x => 229, y => 250),
  (x => 230, y => 250),
  (x => 231, y => 250),
  (x => 237, y => 250),
  (x => 238, y => 250),
  (x => 239, y => 250),
  (x => 240, y => 250),
  (x => 241, y => 250),
  (x => 242, y => 250),
  (x => 246, y => 250),
  (x => 247, y => 250),
  (x => 248, y => 250),
  (x => 258, y => 250),
  (x => 259, y => 250),
  (x => 260, y => 250),
  (x => 261, y => 250),
  (x => 273, y => 250),
  (x => 274, y => 250),
  (x => 275, y => 250),
  (x => 276, y => 250),
  (x => 277, y => 250),
  (x => 278, y => 250),
  (x => 279, y => 250),
  (x => 280, y => 250),
  (x => 281, y => 250),
  (x => 288, y => 250),
  (x => 289, y => 250),
  (x => 290, y => 250),
  (x => 315, y => 250),
  (x => 316, y => 250),
  (x => 317, y => 250),
  (x => 339, y => 250),
  (x => 340, y => 250),
  (x => 341, y => 250),
  (x => 342, y => 250),
  (x => 343, y => 250),
  (x => 353, y => 250),
  (x => 354, y => 250),
  (x => 355, y => 250),
  (x => 356, y => 250),
  (x => 357, y => 250),
  (x => 367, y => 250),
  (x => 368, y => 250),
  (x => 369, y => 250),
  (x => 370, y => 250),
  (x => 376, y => 250),
  (x => 377, y => 250),
  (x => 378, y => 250),
  (x => 379, y => 250),
  (x => 387, y => 250),
  (x => 388, y => 250),
  (x => 389, y => 250),
  (x => 394, y => 250),
  (x => 395, y => 250),
  (x => 396, y => 250),
  (x => 397, y => 250),
  (x => 398, y => 250),
  (x => 399, y => 250),
  (x => 400, y => 250),
  (x => 401, y => 250),
  (x => 402, y => 250),
  (x => 209, y => 251),
  (x => 210, y => 251),
  (x => 211, y => 251),
  (x => 212, y => 251),
  (x => 228, y => 251),
  (x => 229, y => 251),
  (x => 230, y => 251),
  (x => 231, y => 251),
  (x => 238, y => 251),
  (x => 239, y => 251),
  (x => 240, y => 251),
  (x => 241, y => 251),
  (x => 246, y => 251),
  (x => 247, y => 251),
  (x => 248, y => 251),
  (x => 258, y => 251),
  (x => 259, y => 251),
  (x => 260, y => 251),
  (x => 261, y => 251),
  (x => 275, y => 251),
  (x => 276, y => 251),
  (x => 277, y => 251),
  (x => 278, y => 251),
  (x => 279, y => 251),
  (x => 280, y => 251),
  (x => 288, y => 251),
  (x => 289, y => 251),
  (x => 290, y => 251),
  (x => 291, y => 251),
  (x => 315, y => 251),
  (x => 316, y => 251),
  (x => 317, y => 251),
  (x => 340, y => 251),
  (x => 341, y => 251),
  (x => 342, y => 251),
  (x => 343, y => 251),
  (x => 353, y => 251),
  (x => 354, y => 251),
  (x => 355, y => 251),
  (x => 356, y => 251),
  (x => 357, y => 251),
  (x => 367, y => 251),
  (x => 368, y => 251),
  (x => 369, y => 251),
  (x => 370, y => 251),
  (x => 376, y => 251),
  (x => 377, y => 251),
  (x => 378, y => 251),
  (x => 379, y => 251),
  (x => 387, y => 251),
  (x => 388, y => 251),
  (x => 389, y => 251),
  (x => 395, y => 251),
  (x => 396, y => 251),
  (x => 397, y => 251),
  (x => 398, y => 251),
  (x => 399, y => 251),
  (x => 400, y => 251),
  (x => 401, y => 251),
  (x => 258, y => 252),
  (x => 259, y => 252),
  (x => 260, y => 252),
  (x => 261, y => 252),
  (x => 258, y => 253),
  (x => 259, y => 253),
  (x => 260, y => 253),
  (x => 258, y => 254),
  (x => 259, y => 254),
  (x => 260, y => 254),
  (x => 258, y => 255),
  (x => 259, y => 255),
  (x => 260, y => 255),
  (x => 257, y => 256),
  (x => 258, y => 256),
  (x => 259, y => 256),
  (x => 256, y => 257),
  (x => 257, y => 257),
  (x => 258, y => 257),
  (x => 259, y => 257),
  (x => 253, y => 258),
  (x => 254, y => 258),
  (x => 255, y => 258),
  (x => 256, y => 258),
  (x => 257, y => 258),
  (x => 258, y => 258),
  (x => 259, y => 258),
  (x => 253, y => 259),
  (x => 254, y => 259),
  (x => 255, y => 259),
  (x => 256, y => 259),
  (x => 257, y => 259),
  (x => 258, y => 259),
  (x => 253, y => 260),
  (x => 254, y => 260),
  (x => 255, y => 260),
  (x => 256, y => 260),
  (x => 257, y => 260),
  (x => 254, y => 261),
  (x => 255, y => 261)
);
constant p2_end_screen: CoordPairArray(0 to 6614) := (
  (x => 177, y => 128),
  (x => 178, y => 128),
  (x => 179, y => 128),
  (x => 180, y => 128),
  (x => 181, y => 128),
  (x => 182, y => 128),
  (x => 183, y => 128),
  (x => 184, y => 128),
  (x => 185, y => 128),
  (x => 186, y => 128),
  (x => 187, y => 128),
  (x => 188, y => 128),
  (x => 337, y => 128),
  (x => 338, y => 128),
  (x => 339, y => 128),
  (x => 340, y => 128),
  (x => 341, y => 128),
  (x => 342, y => 128),
  (x => 343, y => 128),
  (x => 344, y => 128),
  (x => 345, y => 128),
  (x => 175, y => 129),
  (x => 176, y => 129),
  (x => 177, y => 129),
  (x => 178, y => 129),
  (x => 179, y => 129),
  (x => 180, y => 129),
  (x => 181, y => 129),
  (x => 182, y => 129),
  (x => 183, y => 129),
  (x => 184, y => 129),
  (x => 185, y => 129),
  (x => 186, y => 129),
  (x => 187, y => 129),
  (x => 188, y => 129),
  (x => 189, y => 129),
  (x => 190, y => 129),
  (x => 191, y => 129),
  (x => 334, y => 129),
  (x => 335, y => 129),
  (x => 336, y => 129),
  (x => 337, y => 129),
  (x => 338, y => 129),
  (x => 339, y => 129),
  (x => 340, y => 129),
  (x => 341, y => 129),
  (x => 342, y => 129),
  (x => 343, y => 129),
  (x => 344, y => 129),
  (x => 345, y => 129),
  (x => 346, y => 129),
  (x => 347, y => 129),
  (x => 173, y => 130),
  (x => 174, y => 130),
  (x => 175, y => 130),
  (x => 176, y => 130),
  (x => 177, y => 130),
  (x => 178, y => 130),
  (x => 179, y => 130),
  (x => 180, y => 130),
  (x => 181, y => 130),
  (x => 182, y => 130),
  (x => 183, y => 130),
  (x => 184, y => 130),
  (x => 185, y => 130),
  (x => 186, y => 130),
  (x => 187, y => 130),
  (x => 188, y => 130),
  (x => 189, y => 130),
  (x => 190, y => 130),
  (x => 191, y => 130),
  (x => 333, y => 130),
  (x => 334, y => 130),
  (x => 335, y => 130),
  (x => 336, y => 130),
  (x => 337, y => 130),
  (x => 338, y => 130),
  (x => 339, y => 130),
  (x => 340, y => 130),
  (x => 341, y => 130),
  (x => 342, y => 130),
  (x => 343, y => 130),
  (x => 344, y => 130),
  (x => 345, y => 130),
  (x => 346, y => 130),
  (x => 347, y => 130),
  (x => 348, y => 130),
  (x => 349, y => 130),
  (x => 171, y => 131),
  (x => 172, y => 131),
  (x => 173, y => 131),
  (x => 174, y => 131),
  (x => 175, y => 131),
  (x => 176, y => 131),
  (x => 177, y => 131),
  (x => 178, y => 131),
  (x => 179, y => 131),
  (x => 180, y => 131),
  (x => 181, y => 131),
  (x => 182, y => 131),
  (x => 183, y => 131),
  (x => 184, y => 131),
  (x => 185, y => 131),
  (x => 186, y => 131),
  (x => 187, y => 131),
  (x => 188, y => 131),
  (x => 189, y => 131),
  (x => 190, y => 131),
  (x => 191, y => 131),
  (x => 331, y => 131),
  (x => 332, y => 131),
  (x => 333, y => 131),
  (x => 334, y => 131),
  (x => 335, y => 131),
  (x => 336, y => 131),
  (x => 337, y => 131),
  (x => 338, y => 131),
  (x => 339, y => 131),
  (x => 340, y => 131),
  (x => 341, y => 131),
  (x => 342, y => 131),
  (x => 343, y => 131),
  (x => 344, y => 131),
  (x => 345, y => 131),
  (x => 346, y => 131),
  (x => 347, y => 131),
  (x => 348, y => 131),
  (x => 349, y => 131),
  (x => 350, y => 131),
  (x => 170, y => 132),
  (x => 171, y => 132),
  (x => 172, y => 132),
  (x => 173, y => 132),
  (x => 174, y => 132),
  (x => 175, y => 132),
  (x => 176, y => 132),
  (x => 177, y => 132),
  (x => 178, y => 132),
  (x => 179, y => 132),
  (x => 180, y => 132),
  (x => 181, y => 132),
  (x => 182, y => 132),
  (x => 183, y => 132),
  (x => 184, y => 132),
  (x => 185, y => 132),
  (x => 186, y => 132),
  (x => 187, y => 132),
  (x => 188, y => 132),
  (x => 189, y => 132),
  (x => 190, y => 132),
  (x => 191, y => 132),
  (x => 330, y => 132),
  (x => 331, y => 132),
  (x => 332, y => 132),
  (x => 333, y => 132),
  (x => 334, y => 132),
  (x => 335, y => 132),
  (x => 336, y => 132),
  (x => 337, y => 132),
  (x => 338, y => 132),
  (x => 339, y => 132),
  (x => 340, y => 132),
  (x => 341, y => 132),
  (x => 342, y => 132),
  (x => 343, y => 132),
  (x => 344, y => 132),
  (x => 345, y => 132),
  (x => 346, y => 132),
  (x => 347, y => 132),
  (x => 348, y => 132),
  (x => 349, y => 132),
  (x => 350, y => 132),
  (x => 351, y => 132),
  (x => 169, y => 133),
  (x => 170, y => 133),
  (x => 171, y => 133),
  (x => 172, y => 133),
  (x => 173, y => 133),
  (x => 174, y => 133),
  (x => 175, y => 133),
  (x => 176, y => 133),
  (x => 177, y => 133),
  (x => 178, y => 133),
  (x => 179, y => 133),
  (x => 180, y => 133),
  (x => 181, y => 133),
  (x => 182, y => 133),
  (x => 183, y => 133),
  (x => 184, y => 133),
  (x => 185, y => 133),
  (x => 186, y => 133),
  (x => 187, y => 133),
  (x => 188, y => 133),
  (x => 189, y => 133),
  (x => 190, y => 133),
  (x => 191, y => 133),
  (x => 329, y => 133),
  (x => 330, y => 133),
  (x => 331, y => 133),
  (x => 332, y => 133),
  (x => 333, y => 133),
  (x => 334, y => 133),
  (x => 335, y => 133),
  (x => 336, y => 133),
  (x => 337, y => 133),
  (x => 338, y => 133),
  (x => 339, y => 133),
  (x => 340, y => 133),
  (x => 341, y => 133),
  (x => 342, y => 133),
  (x => 343, y => 133),
  (x => 344, y => 133),
  (x => 345, y => 133),
  (x => 346, y => 133),
  (x => 347, y => 133),
  (x => 348, y => 133),
  (x => 349, y => 133),
  (x => 350, y => 133),
  (x => 351, y => 133),
  (x => 352, y => 133),
  (x => 168, y => 134),
  (x => 169, y => 134),
  (x => 170, y => 134),
  (x => 171, y => 134),
  (x => 172, y => 134),
  (x => 173, y => 134),
  (x => 174, y => 134),
  (x => 175, y => 134),
  (x => 176, y => 134),
  (x => 177, y => 134),
  (x => 178, y => 134),
  (x => 179, y => 134),
  (x => 180, y => 134),
  (x => 181, y => 134),
  (x => 182, y => 134),
  (x => 183, y => 134),
  (x => 184, y => 134),
  (x => 185, y => 134),
  (x => 186, y => 134),
  (x => 187, y => 134),
  (x => 188, y => 134),
  (x => 189, y => 134),
  (x => 190, y => 134),
  (x => 191, y => 134),
  (x => 329, y => 134),
  (x => 330, y => 134),
  (x => 331, y => 134),
  (x => 332, y => 134),
  (x => 333, y => 134),
  (x => 334, y => 134),
  (x => 335, y => 134),
  (x => 336, y => 134),
  (x => 337, y => 134),
  (x => 338, y => 134),
  (x => 339, y => 134),
  (x => 340, y => 134),
  (x => 341, y => 134),
  (x => 342, y => 134),
  (x => 343, y => 134),
  (x => 344, y => 134),
  (x => 345, y => 134),
  (x => 346, y => 134),
  (x => 347, y => 134),
  (x => 348, y => 134),
  (x => 349, y => 134),
  (x => 350, y => 134),
  (x => 351, y => 134),
  (x => 352, y => 134),
  (x => 353, y => 134),
  (x => 167, y => 135),
  (x => 168, y => 135),
  (x => 169, y => 135),
  (x => 170, y => 135),
  (x => 171, y => 135),
  (x => 172, y => 135),
  (x => 173, y => 135),
  (x => 174, y => 135),
  (x => 175, y => 135),
  (x => 176, y => 135),
  (x => 177, y => 135),
  (x => 178, y => 135),
  (x => 179, y => 135),
  (x => 180, y => 135),
  (x => 181, y => 135),
  (x => 182, y => 135),
  (x => 183, y => 135),
  (x => 184, y => 135),
  (x => 185, y => 135),
  (x => 186, y => 135),
  (x => 187, y => 135),
  (x => 188, y => 135),
  (x => 189, y => 135),
  (x => 190, y => 135),
  (x => 191, y => 135),
  (x => 328, y => 135),
  (x => 329, y => 135),
  (x => 330, y => 135),
  (x => 331, y => 135),
  (x => 332, y => 135),
  (x => 333, y => 135),
  (x => 334, y => 135),
  (x => 335, y => 135),
  (x => 336, y => 135),
  (x => 337, y => 135),
  (x => 338, y => 135),
  (x => 339, y => 135),
  (x => 340, y => 135),
  (x => 341, y => 135),
  (x => 342, y => 135),
  (x => 343, y => 135),
  (x => 344, y => 135),
  (x => 345, y => 135),
  (x => 346, y => 135),
  (x => 347, y => 135),
  (x => 348, y => 135),
  (x => 349, y => 135),
  (x => 350, y => 135),
  (x => 351, y => 135),
  (x => 352, y => 135),
  (x => 353, y => 135),
  (x => 354, y => 135),
  (x => 167, y => 136),
  (x => 168, y => 136),
  (x => 169, y => 136),
  (x => 170, y => 136),
  (x => 171, y => 136),
  (x => 172, y => 136),
  (x => 173, y => 136),
  (x => 174, y => 136),
  (x => 175, y => 136),
  (x => 176, y => 136),
  (x => 177, y => 136),
  (x => 178, y => 136),
  (x => 188, y => 136),
  (x => 189, y => 136),
  (x => 190, y => 136),
  (x => 191, y => 136),
  (x => 327, y => 136),
  (x => 328, y => 136),
  (x => 329, y => 136),
  (x => 330, y => 136),
  (x => 331, y => 136),
  (x => 332, y => 136),
  (x => 333, y => 136),
  (x => 334, y => 136),
  (x => 335, y => 136),
  (x => 336, y => 136),
  (x => 337, y => 136),
  (x => 338, y => 136),
  (x => 344, y => 136),
  (x => 345, y => 136),
  (x => 346, y => 136),
  (x => 347, y => 136),
  (x => 348, y => 136),
  (x => 349, y => 136),
  (x => 350, y => 136),
  (x => 351, y => 136),
  (x => 352, y => 136),
  (x => 353, y => 136),
  (x => 354, y => 136),
  (x => 166, y => 137),
  (x => 167, y => 137),
  (x => 168, y => 137),
  (x => 169, y => 137),
  (x => 170, y => 137),
  (x => 171, y => 137),
  (x => 172, y => 137),
  (x => 173, y => 137),
  (x => 174, y => 137),
  (x => 175, y => 137),
  (x => 176, y => 137),
  (x => 190, y => 137),
  (x => 191, y => 137),
  (x => 327, y => 137),
  (x => 328, y => 137),
  (x => 329, y => 137),
  (x => 330, y => 137),
  (x => 331, y => 137),
  (x => 332, y => 137),
  (x => 333, y => 137),
  (x => 334, y => 137),
  (x => 335, y => 137),
  (x => 336, y => 137),
  (x => 346, y => 137),
  (x => 347, y => 137),
  (x => 348, y => 137),
  (x => 349, y => 137),
  (x => 350, y => 137),
  (x => 351, y => 137),
  (x => 352, y => 137),
  (x => 353, y => 137),
  (x => 354, y => 137),
  (x => 355, y => 137),
  (x => 166, y => 138),
  (x => 167, y => 138),
  (x => 168, y => 138),
  (x => 169, y => 138),
  (x => 170, y => 138),
  (x => 171, y => 138),
  (x => 172, y => 138),
  (x => 173, y => 138),
  (x => 174, y => 138),
  (x => 326, y => 138),
  (x => 327, y => 138),
  (x => 328, y => 138),
  (x => 329, y => 138),
  (x => 330, y => 138),
  (x => 331, y => 138),
  (x => 332, y => 138),
  (x => 333, y => 138),
  (x => 334, y => 138),
  (x => 347, y => 138),
  (x => 348, y => 138),
  (x => 349, y => 138),
  (x => 350, y => 138),
  (x => 351, y => 138),
  (x => 352, y => 138),
  (x => 353, y => 138),
  (x => 354, y => 138),
  (x => 355, y => 138),
  (x => 165, y => 139),
  (x => 166, y => 139),
  (x => 167, y => 139),
  (x => 168, y => 139),
  (x => 169, y => 139),
  (x => 170, y => 139),
  (x => 171, y => 139),
  (x => 172, y => 139),
  (x => 173, y => 139),
  (x => 326, y => 139),
  (x => 327, y => 139),
  (x => 328, y => 139),
  (x => 329, y => 139),
  (x => 330, y => 139),
  (x => 331, y => 139),
  (x => 332, y => 139),
  (x => 333, y => 139),
  (x => 334, y => 139),
  (x => 348, y => 139),
  (x => 349, y => 139),
  (x => 350, y => 139),
  (x => 351, y => 139),
  (x => 352, y => 139),
  (x => 353, y => 139),
  (x => 354, y => 139),
  (x => 355, y => 139),
  (x => 356, y => 139),
  (x => 165, y => 140),
  (x => 166, y => 140),
  (x => 167, y => 140),
  (x => 168, y => 140),
  (x => 169, y => 140),
  (x => 170, y => 140),
  (x => 171, y => 140),
  (x => 172, y => 140),
  (x => 325, y => 140),
  (x => 326, y => 140),
  (x => 327, y => 140),
  (x => 328, y => 140),
  (x => 329, y => 140),
  (x => 330, y => 140),
  (x => 331, y => 140),
  (x => 332, y => 140),
  (x => 333, y => 140),
  (x => 348, y => 140),
  (x => 349, y => 140),
  (x => 350, y => 140),
  (x => 351, y => 140),
  (x => 352, y => 140),
  (x => 353, y => 140),
  (x => 354, y => 140),
  (x => 355, y => 140),
  (x => 356, y => 140),
  (x => 164, y => 141),
  (x => 165, y => 141),
  (x => 166, y => 141),
  (x => 167, y => 141),
  (x => 168, y => 141),
  (x => 169, y => 141),
  (x => 170, y => 141),
  (x => 171, y => 141),
  (x => 172, y => 141),
  (x => 325, y => 141),
  (x => 326, y => 141),
  (x => 327, y => 141),
  (x => 328, y => 141),
  (x => 329, y => 141),
  (x => 330, y => 141),
  (x => 331, y => 141),
  (x => 332, y => 141),
  (x => 349, y => 141),
  (x => 350, y => 141),
  (x => 351, y => 141),
  (x => 352, y => 141),
  (x => 353, y => 141),
  (x => 354, y => 141),
  (x => 355, y => 141),
  (x => 356, y => 141),
  (x => 164, y => 142),
  (x => 165, y => 142),
  (x => 166, y => 142),
  (x => 167, y => 142),
  (x => 168, y => 142),
  (x => 169, y => 142),
  (x => 170, y => 142),
  (x => 171, y => 142),
  (x => 210, y => 142),
  (x => 211, y => 142),
  (x => 212, y => 142),
  (x => 213, y => 142),
  (x => 214, y => 142),
  (x => 246, y => 142),
  (x => 247, y => 142),
  (x => 248, y => 142),
  (x => 263, y => 142),
  (x => 264, y => 142),
  (x => 265, y => 142),
  (x => 290, y => 142),
  (x => 291, y => 142),
  (x => 292, y => 142),
  (x => 293, y => 142),
  (x => 325, y => 142),
  (x => 326, y => 142),
  (x => 327, y => 142),
  (x => 328, y => 142),
  (x => 329, y => 142),
  (x => 330, y => 142),
  (x => 331, y => 142),
  (x => 332, y => 142),
  (x => 350, y => 142),
  (x => 351, y => 142),
  (x => 352, y => 142),
  (x => 353, y => 142),
  (x => 354, y => 142),
  (x => 355, y => 142),
  (x => 356, y => 142),
  (x => 357, y => 142),
  (x => 404, y => 142),
  (x => 405, y => 142),
  (x => 406, y => 142),
  (x => 407, y => 142),
  (x => 438, y => 142),
  (x => 439, y => 142),
  (x => 164, y => 143),
  (x => 165, y => 143),
  (x => 166, y => 143),
  (x => 167, y => 143),
  (x => 168, y => 143),
  (x => 169, y => 143),
  (x => 170, y => 143),
  (x => 171, y => 143),
  (x => 206, y => 143),
  (x => 207, y => 143),
  (x => 208, y => 143),
  (x => 209, y => 143),
  (x => 210, y => 143),
  (x => 211, y => 143),
  (x => 212, y => 143),
  (x => 213, y => 143),
  (x => 214, y => 143),
  (x => 215, y => 143),
  (x => 216, y => 143),
  (x => 217, y => 143),
  (x => 231, y => 143),
  (x => 232, y => 143),
  (x => 233, y => 143),
  (x => 234, y => 143),
  (x => 235, y => 143),
  (x => 236, y => 143),
  (x => 237, y => 143),
  (x => 243, y => 143),
  (x => 244, y => 143),
  (x => 245, y => 143),
  (x => 246, y => 143),
  (x => 247, y => 143),
  (x => 248, y => 143),
  (x => 249, y => 143),
  (x => 250, y => 143),
  (x => 251, y => 143),
  (x => 260, y => 143),
  (x => 261, y => 143),
  (x => 262, y => 143),
  (x => 263, y => 143),
  (x => 264, y => 143),
  (x => 265, y => 143),
  (x => 266, y => 143),
  (x => 267, y => 143),
  (x => 268, y => 143),
  (x => 287, y => 143),
  (x => 288, y => 143),
  (x => 289, y => 143),
  (x => 290, y => 143),
  (x => 291, y => 143),
  (x => 292, y => 143),
  (x => 293, y => 143),
  (x => 294, y => 143),
  (x => 295, y => 143),
  (x => 296, y => 143),
  (x => 324, y => 143),
  (x => 325, y => 143),
  (x => 326, y => 143),
  (x => 327, y => 143),
  (x => 328, y => 143),
  (x => 329, y => 143),
  (x => 330, y => 143),
  (x => 331, y => 143),
  (x => 350, y => 143),
  (x => 351, y => 143),
  (x => 352, y => 143),
  (x => 353, y => 143),
  (x => 354, y => 143),
  (x => 355, y => 143),
  (x => 356, y => 143),
  (x => 357, y => 143),
  (x => 362, y => 143),
  (x => 363, y => 143),
  (x => 364, y => 143),
  (x => 365, y => 143),
  (x => 366, y => 143),
  (x => 367, y => 143),
  (x => 368, y => 143),
  (x => 369, y => 143),
  (x => 382, y => 143),
  (x => 383, y => 143),
  (x => 384, y => 143),
  (x => 385, y => 143),
  (x => 386, y => 143),
  (x => 387, y => 143),
  (x => 388, y => 143),
  (x => 389, y => 143),
  (x => 401, y => 143),
  (x => 402, y => 143),
  (x => 403, y => 143),
  (x => 404, y => 143),
  (x => 405, y => 143),
  (x => 406, y => 143),
  (x => 407, y => 143),
  (x => 408, y => 143),
  (x => 409, y => 143),
  (x => 410, y => 143),
  (x => 424, y => 143),
  (x => 425, y => 143),
  (x => 426, y => 143),
  (x => 427, y => 143),
  (x => 428, y => 143),
  (x => 429, y => 143),
  (x => 430, y => 143),
  (x => 436, y => 143),
  (x => 437, y => 143),
  (x => 438, y => 143),
  (x => 439, y => 143),
  (x => 163, y => 144),
  (x => 164, y => 144),
  (x => 165, y => 144),
  (x => 166, y => 144),
  (x => 167, y => 144),
  (x => 168, y => 144),
  (x => 169, y => 144),
  (x => 170, y => 144),
  (x => 204, y => 144),
  (x => 205, y => 144),
  (x => 206, y => 144),
  (x => 207, y => 144),
  (x => 208, y => 144),
  (x => 209, y => 144),
  (x => 210, y => 144),
  (x => 211, y => 144),
  (x => 212, y => 144),
  (x => 213, y => 144),
  (x => 214, y => 144),
  (x => 215, y => 144),
  (x => 216, y => 144),
  (x => 217, y => 144),
  (x => 218, y => 144),
  (x => 231, y => 144),
  (x => 232, y => 144),
  (x => 233, y => 144),
  (x => 234, y => 144),
  (x => 235, y => 144),
  (x => 236, y => 144),
  (x => 237, y => 144),
  (x => 242, y => 144),
  (x => 243, y => 144),
  (x => 244, y => 144),
  (x => 245, y => 144),
  (x => 246, y => 144),
  (x => 247, y => 144),
  (x => 248, y => 144),
  (x => 249, y => 144),
  (x => 250, y => 144),
  (x => 251, y => 144),
  (x => 252, y => 144),
  (x => 259, y => 144),
  (x => 260, y => 144),
  (x => 261, y => 144),
  (x => 262, y => 144),
  (x => 263, y => 144),
  (x => 264, y => 144),
  (x => 265, y => 144),
  (x => 266, y => 144),
  (x => 267, y => 144),
  (x => 268, y => 144),
  (x => 269, y => 144),
  (x => 285, y => 144),
  (x => 286, y => 144),
  (x => 287, y => 144),
  (x => 288, y => 144),
  (x => 289, y => 144),
  (x => 290, y => 144),
  (x => 291, y => 144),
  (x => 292, y => 144),
  (x => 293, y => 144),
  (x => 294, y => 144),
  (x => 295, y => 144),
  (x => 296, y => 144),
  (x => 297, y => 144),
  (x => 324, y => 144),
  (x => 325, y => 144),
  (x => 326, y => 144),
  (x => 327, y => 144),
  (x => 328, y => 144),
  (x => 329, y => 144),
  (x => 330, y => 144),
  (x => 331, y => 144),
  (x => 350, y => 144),
  (x => 351, y => 144),
  (x => 352, y => 144),
  (x => 353, y => 144),
  (x => 354, y => 144),
  (x => 355, y => 144),
  (x => 356, y => 144),
  (x => 357, y => 144),
  (x => 363, y => 144),
  (x => 364, y => 144),
  (x => 365, y => 144),
  (x => 366, y => 144),
  (x => 367, y => 144),
  (x => 368, y => 144),
  (x => 369, y => 144),
  (x => 382, y => 144),
  (x => 383, y => 144),
  (x => 384, y => 144),
  (x => 385, y => 144),
  (x => 386, y => 144),
  (x => 387, y => 144),
  (x => 388, y => 144),
  (x => 400, y => 144),
  (x => 401, y => 144),
  (x => 402, y => 144),
  (x => 403, y => 144),
  (x => 404, y => 144),
  (x => 405, y => 144),
  (x => 406, y => 144),
  (x => 407, y => 144),
  (x => 408, y => 144),
  (x => 409, y => 144),
  (x => 410, y => 144),
  (x => 411, y => 144),
  (x => 412, y => 144),
  (x => 424, y => 144),
  (x => 425, y => 144),
  (x => 426, y => 144),
  (x => 427, y => 144),
  (x => 428, y => 144),
  (x => 429, y => 144),
  (x => 430, y => 144),
  (x => 435, y => 144),
  (x => 436, y => 144),
  (x => 437, y => 144),
  (x => 438, y => 144),
  (x => 439, y => 144),
  (x => 163, y => 145),
  (x => 164, y => 145),
  (x => 165, y => 145),
  (x => 166, y => 145),
  (x => 167, y => 145),
  (x => 168, y => 145),
  (x => 169, y => 145),
  (x => 170, y => 145),
  (x => 203, y => 145),
  (x => 204, y => 145),
  (x => 205, y => 145),
  (x => 206, y => 145),
  (x => 207, y => 145),
  (x => 208, y => 145),
  (x => 209, y => 145),
  (x => 210, y => 145),
  (x => 211, y => 145),
  (x => 212, y => 145),
  (x => 213, y => 145),
  (x => 214, y => 145),
  (x => 215, y => 145),
  (x => 216, y => 145),
  (x => 217, y => 145),
  (x => 218, y => 145),
  (x => 219, y => 145),
  (x => 231, y => 145),
  (x => 232, y => 145),
  (x => 233, y => 145),
  (x => 234, y => 145),
  (x => 235, y => 145),
  (x => 236, y => 145),
  (x => 237, y => 145),
  (x => 241, y => 145),
  (x => 242, y => 145),
  (x => 243, y => 145),
  (x => 244, y => 145),
  (x => 245, y => 145),
  (x => 246, y => 145),
  (x => 247, y => 145),
  (x => 248, y => 145),
  (x => 249, y => 145),
  (x => 250, y => 145),
  (x => 251, y => 145),
  (x => 252, y => 145),
  (x => 258, y => 145),
  (x => 259, y => 145),
  (x => 260, y => 145),
  (x => 261, y => 145),
  (x => 262, y => 145),
  (x => 263, y => 145),
  (x => 264, y => 145),
  (x => 265, y => 145),
  (x => 266, y => 145),
  (x => 267, y => 145),
  (x => 268, y => 145),
  (x => 269, y => 145),
  (x => 284, y => 145),
  (x => 285, y => 145),
  (x => 286, y => 145),
  (x => 287, y => 145),
  (x => 288, y => 145),
  (x => 289, y => 145),
  (x => 290, y => 145),
  (x => 291, y => 145),
  (x => 292, y => 145),
  (x => 293, y => 145),
  (x => 294, y => 145),
  (x => 295, y => 145),
  (x => 296, y => 145),
  (x => 297, y => 145),
  (x => 298, y => 145),
  (x => 324, y => 145),
  (x => 325, y => 145),
  (x => 326, y => 145),
  (x => 327, y => 145),
  (x => 328, y => 145),
  (x => 329, y => 145),
  (x => 330, y => 145),
  (x => 331, y => 145),
  (x => 350, y => 145),
  (x => 351, y => 145),
  (x => 352, y => 145),
  (x => 353, y => 145),
  (x => 354, y => 145),
  (x => 355, y => 145),
  (x => 356, y => 145),
  (x => 357, y => 145),
  (x => 363, y => 145),
  (x => 364, y => 145),
  (x => 365, y => 145),
  (x => 366, y => 145),
  (x => 367, y => 145),
  (x => 368, y => 145),
  (x => 369, y => 145),
  (x => 382, y => 145),
  (x => 383, y => 145),
  (x => 384, y => 145),
  (x => 385, y => 145),
  (x => 386, y => 145),
  (x => 387, y => 145),
  (x => 388, y => 145),
  (x => 399, y => 145),
  (x => 400, y => 145),
  (x => 401, y => 145),
  (x => 402, y => 145),
  (x => 403, y => 145),
  (x => 404, y => 145),
  (x => 405, y => 145),
  (x => 406, y => 145),
  (x => 407, y => 145),
  (x => 408, y => 145),
  (x => 409, y => 145),
  (x => 410, y => 145),
  (x => 411, y => 145),
  (x => 412, y => 145),
  (x => 413, y => 145),
  (x => 424, y => 145),
  (x => 425, y => 145),
  (x => 426, y => 145),
  (x => 427, y => 145),
  (x => 428, y => 145),
  (x => 429, y => 145),
  (x => 430, y => 145),
  (x => 434, y => 145),
  (x => 435, y => 145),
  (x => 436, y => 145),
  (x => 437, y => 145),
  (x => 438, y => 145),
  (x => 439, y => 145),
  (x => 163, y => 146),
  (x => 164, y => 146),
  (x => 165, y => 146),
  (x => 166, y => 146),
  (x => 167, y => 146),
  (x => 168, y => 146),
  (x => 169, y => 146),
  (x => 170, y => 146),
  (x => 203, y => 146),
  (x => 204, y => 146),
  (x => 205, y => 146),
  (x => 206, y => 146),
  (x => 207, y => 146),
  (x => 208, y => 146),
  (x => 209, y => 146),
  (x => 210, y => 146),
  (x => 211, y => 146),
  (x => 212, y => 146),
  (x => 213, y => 146),
  (x => 214, y => 146),
  (x => 215, y => 146),
  (x => 216, y => 146),
  (x => 217, y => 146),
  (x => 218, y => 146),
  (x => 219, y => 146),
  (x => 220, y => 146),
  (x => 231, y => 146),
  (x => 232, y => 146),
  (x => 233, y => 146),
  (x => 234, y => 146),
  (x => 235, y => 146),
  (x => 236, y => 146),
  (x => 237, y => 146),
  (x => 240, y => 146),
  (x => 241, y => 146),
  (x => 242, y => 146),
  (x => 243, y => 146),
  (x => 244, y => 146),
  (x => 245, y => 146),
  (x => 246, y => 146),
  (x => 247, y => 146),
  (x => 248, y => 146),
  (x => 249, y => 146),
  (x => 250, y => 146),
  (x => 251, y => 146),
  (x => 252, y => 146),
  (x => 253, y => 146),
  (x => 257, y => 146),
  (x => 258, y => 146),
  (x => 259, y => 146),
  (x => 260, y => 146),
  (x => 261, y => 146),
  (x => 262, y => 146),
  (x => 263, y => 146),
  (x => 264, y => 146),
  (x => 265, y => 146),
  (x => 266, y => 146),
  (x => 267, y => 146),
  (x => 268, y => 146),
  (x => 269, y => 146),
  (x => 270, y => 146),
  (x => 283, y => 146),
  (x => 284, y => 146),
  (x => 285, y => 146),
  (x => 286, y => 146),
  (x => 287, y => 146),
  (x => 288, y => 146),
  (x => 289, y => 146),
  (x => 290, y => 146),
  (x => 291, y => 146),
  (x => 292, y => 146),
  (x => 293, y => 146),
  (x => 294, y => 146),
  (x => 295, y => 146),
  (x => 296, y => 146),
  (x => 297, y => 146),
  (x => 298, y => 146),
  (x => 299, y => 146),
  (x => 324, y => 146),
  (x => 325, y => 146),
  (x => 326, y => 146),
  (x => 327, y => 146),
  (x => 328, y => 146),
  (x => 329, y => 146),
  (x => 330, y => 146),
  (x => 351, y => 146),
  (x => 352, y => 146),
  (x => 353, y => 146),
  (x => 354, y => 146),
  (x => 355, y => 146),
  (x => 356, y => 146),
  (x => 357, y => 146),
  (x => 363, y => 146),
  (x => 364, y => 146),
  (x => 365, y => 146),
  (x => 366, y => 146),
  (x => 367, y => 146),
  (x => 368, y => 146),
  (x => 369, y => 146),
  (x => 370, y => 146),
  (x => 382, y => 146),
  (x => 383, y => 146),
  (x => 384, y => 146),
  (x => 385, y => 146),
  (x => 386, y => 146),
  (x => 387, y => 146),
  (x => 388, y => 146),
  (x => 398, y => 146),
  (x => 399, y => 146),
  (x => 400, y => 146),
  (x => 401, y => 146),
  (x => 402, y => 146),
  (x => 403, y => 146),
  (x => 404, y => 146),
  (x => 405, y => 146),
  (x => 406, y => 146),
  (x => 407, y => 146),
  (x => 408, y => 146),
  (x => 409, y => 146),
  (x => 410, y => 146),
  (x => 411, y => 146),
  (x => 412, y => 146),
  (x => 413, y => 146),
  (x => 414, y => 146),
  (x => 424, y => 146),
  (x => 425, y => 146),
  (x => 426, y => 146),
  (x => 427, y => 146),
  (x => 428, y => 146),
  (x => 429, y => 146),
  (x => 430, y => 146),
  (x => 434, y => 146),
  (x => 435, y => 146),
  (x => 436, y => 146),
  (x => 437, y => 146),
  (x => 438, y => 146),
  (x => 439, y => 146),
  (x => 163, y => 147),
  (x => 164, y => 147),
  (x => 165, y => 147),
  (x => 166, y => 147),
  (x => 167, y => 147),
  (x => 168, y => 147),
  (x => 169, y => 147),
  (x => 203, y => 147),
  (x => 204, y => 147),
  (x => 205, y => 147),
  (x => 206, y => 147),
  (x => 207, y => 147),
  (x => 208, y => 147),
  (x => 209, y => 147),
  (x => 210, y => 147),
  (x => 211, y => 147),
  (x => 212, y => 147),
  (x => 213, y => 147),
  (x => 214, y => 147),
  (x => 215, y => 147),
  (x => 216, y => 147),
  (x => 217, y => 147),
  (x => 218, y => 147),
  (x => 219, y => 147),
  (x => 220, y => 147),
  (x => 231, y => 147),
  (x => 232, y => 147),
  (x => 233, y => 147),
  (x => 234, y => 147),
  (x => 235, y => 147),
  (x => 236, y => 147),
  (x => 237, y => 147),
  (x => 240, y => 147),
  (x => 241, y => 147),
  (x => 242, y => 147),
  (x => 243, y => 147),
  (x => 244, y => 147),
  (x => 245, y => 147),
  (x => 246, y => 147),
  (x => 247, y => 147),
  (x => 248, y => 147),
  (x => 249, y => 147),
  (x => 250, y => 147),
  (x => 251, y => 147),
  (x => 252, y => 147),
  (x => 253, y => 147),
  (x => 257, y => 147),
  (x => 258, y => 147),
  (x => 259, y => 147),
  (x => 260, y => 147),
  (x => 261, y => 147),
  (x => 262, y => 147),
  (x => 263, y => 147),
  (x => 264, y => 147),
  (x => 265, y => 147),
  (x => 266, y => 147),
  (x => 267, y => 147),
  (x => 268, y => 147),
  (x => 269, y => 147),
  (x => 270, y => 147),
  (x => 282, y => 147),
  (x => 283, y => 147),
  (x => 284, y => 147),
  (x => 285, y => 147),
  (x => 286, y => 147),
  (x => 287, y => 147),
  (x => 288, y => 147),
  (x => 289, y => 147),
  (x => 290, y => 147),
  (x => 291, y => 147),
  (x => 292, y => 147),
  (x => 293, y => 147),
  (x => 294, y => 147),
  (x => 295, y => 147),
  (x => 296, y => 147),
  (x => 297, y => 147),
  (x => 298, y => 147),
  (x => 299, y => 147),
  (x => 300, y => 147),
  (x => 324, y => 147),
  (x => 325, y => 147),
  (x => 326, y => 147),
  (x => 327, y => 147),
  (x => 328, y => 147),
  (x => 329, y => 147),
  (x => 330, y => 147),
  (x => 351, y => 147),
  (x => 352, y => 147),
  (x => 353, y => 147),
  (x => 354, y => 147),
  (x => 355, y => 147),
  (x => 356, y => 147),
  (x => 357, y => 147),
  (x => 358, y => 147),
  (x => 364, y => 147),
  (x => 365, y => 147),
  (x => 366, y => 147),
  (x => 367, y => 147),
  (x => 368, y => 147),
  (x => 369, y => 147),
  (x => 370, y => 147),
  (x => 382, y => 147),
  (x => 383, y => 147),
  (x => 384, y => 147),
  (x => 385, y => 147),
  (x => 386, y => 147),
  (x => 387, y => 147),
  (x => 388, y => 147),
  (x => 397, y => 147),
  (x => 398, y => 147),
  (x => 399, y => 147),
  (x => 400, y => 147),
  (x => 401, y => 147),
  (x => 402, y => 147),
  (x => 403, y => 147),
  (x => 404, y => 147),
  (x => 405, y => 147),
  (x => 406, y => 147),
  (x => 407, y => 147),
  (x => 408, y => 147),
  (x => 409, y => 147),
  (x => 410, y => 147),
  (x => 411, y => 147),
  (x => 412, y => 147),
  (x => 413, y => 147),
  (x => 414, y => 147),
  (x => 424, y => 147),
  (x => 425, y => 147),
  (x => 426, y => 147),
  (x => 427, y => 147),
  (x => 428, y => 147),
  (x => 429, y => 147),
  (x => 430, y => 147),
  (x => 433, y => 147),
  (x => 434, y => 147),
  (x => 435, y => 147),
  (x => 436, y => 147),
  (x => 437, y => 147),
  (x => 438, y => 147),
  (x => 439, y => 147),
  (x => 163, y => 148),
  (x => 164, y => 148),
  (x => 165, y => 148),
  (x => 166, y => 148),
  (x => 167, y => 148),
  (x => 168, y => 148),
  (x => 169, y => 148),
  (x => 203, y => 148),
  (x => 204, y => 148),
  (x => 205, y => 148),
  (x => 206, y => 148),
  (x => 207, y => 148),
  (x => 208, y => 148),
  (x => 213, y => 148),
  (x => 214, y => 148),
  (x => 215, y => 148),
  (x => 216, y => 148),
  (x => 217, y => 148),
  (x => 218, y => 148),
  (x => 219, y => 148),
  (x => 220, y => 148),
  (x => 221, y => 148),
  (x => 231, y => 148),
  (x => 232, y => 148),
  (x => 233, y => 148),
  (x => 234, y => 148),
  (x => 235, y => 148),
  (x => 236, y => 148),
  (x => 237, y => 148),
  (x => 239, y => 148),
  (x => 240, y => 148),
  (x => 241, y => 148),
  (x => 242, y => 148),
  (x => 243, y => 148),
  (x => 244, y => 148),
  (x => 245, y => 148),
  (x => 246, y => 148),
  (x => 247, y => 148),
  (x => 248, y => 148),
  (x => 249, y => 148),
  (x => 250, y => 148),
  (x => 251, y => 148),
  (x => 252, y => 148),
  (x => 253, y => 148),
  (x => 254, y => 148),
  (x => 256, y => 148),
  (x => 257, y => 148),
  (x => 258, y => 148),
  (x => 259, y => 148),
  (x => 260, y => 148),
  (x => 261, y => 148),
  (x => 262, y => 148),
  (x => 263, y => 148),
  (x => 264, y => 148),
  (x => 265, y => 148),
  (x => 266, y => 148),
  (x => 267, y => 148),
  (x => 268, y => 148),
  (x => 269, y => 148),
  (x => 270, y => 148),
  (x => 271, y => 148),
  (x => 282, y => 148),
  (x => 283, y => 148),
  (x => 284, y => 148),
  (x => 285, y => 148),
  (x => 286, y => 148),
  (x => 287, y => 148),
  (x => 288, y => 148),
  (x => 289, y => 148),
  (x => 293, y => 148),
  (x => 294, y => 148),
  (x => 295, y => 148),
  (x => 296, y => 148),
  (x => 297, y => 148),
  (x => 298, y => 148),
  (x => 299, y => 148),
  (x => 300, y => 148),
  (x => 324, y => 148),
  (x => 325, y => 148),
  (x => 326, y => 148),
  (x => 327, y => 148),
  (x => 328, y => 148),
  (x => 329, y => 148),
  (x => 330, y => 148),
  (x => 351, y => 148),
  (x => 352, y => 148),
  (x => 353, y => 148),
  (x => 354, y => 148),
  (x => 355, y => 148),
  (x => 356, y => 148),
  (x => 357, y => 148),
  (x => 358, y => 148),
  (x => 364, y => 148),
  (x => 365, y => 148),
  (x => 366, y => 148),
  (x => 367, y => 148),
  (x => 368, y => 148),
  (x => 369, y => 148),
  (x => 370, y => 148),
  (x => 382, y => 148),
  (x => 383, y => 148),
  (x => 384, y => 148),
  (x => 385, y => 148),
  (x => 386, y => 148),
  (x => 387, y => 148),
  (x => 396, y => 148),
  (x => 397, y => 148),
  (x => 398, y => 148),
  (x => 399, y => 148),
  (x => 400, y => 148),
  (x => 401, y => 148),
  (x => 402, y => 148),
  (x => 403, y => 148),
  (x => 404, y => 148),
  (x => 408, y => 148),
  (x => 409, y => 148),
  (x => 410, y => 148),
  (x => 411, y => 148),
  (x => 412, y => 148),
  (x => 413, y => 148),
  (x => 414, y => 148),
  (x => 415, y => 148),
  (x => 424, y => 148),
  (x => 425, y => 148),
  (x => 426, y => 148),
  (x => 427, y => 148),
  (x => 428, y => 148),
  (x => 429, y => 148),
  (x => 430, y => 148),
  (x => 433, y => 148),
  (x => 434, y => 148),
  (x => 435, y => 148),
  (x => 436, y => 148),
  (x => 437, y => 148),
  (x => 438, y => 148),
  (x => 439, y => 148),
  (x => 162, y => 149),
  (x => 163, y => 149),
  (x => 164, y => 149),
  (x => 165, y => 149),
  (x => 166, y => 149),
  (x => 167, y => 149),
  (x => 168, y => 149),
  (x => 169, y => 149),
  (x => 203, y => 149),
  (x => 204, y => 149),
  (x => 205, y => 149),
  (x => 215, y => 149),
  (x => 216, y => 149),
  (x => 217, y => 149),
  (x => 218, y => 149),
  (x => 219, y => 149),
  (x => 220, y => 149),
  (x => 221, y => 149),
  (x => 231, y => 149),
  (x => 232, y => 149),
  (x => 233, y => 149),
  (x => 234, y => 149),
  (x => 235, y => 149),
  (x => 236, y => 149),
  (x => 237, y => 149),
  (x => 238, y => 149),
  (x => 239, y => 149),
  (x => 240, y => 149),
  (x => 241, y => 149),
  (x => 245, y => 149),
  (x => 246, y => 149),
  (x => 247, y => 149),
  (x => 248, y => 149),
  (x => 249, y => 149),
  (x => 250, y => 149),
  (x => 251, y => 149),
  (x => 252, y => 149),
  (x => 253, y => 149),
  (x => 254, y => 149),
  (x => 255, y => 149),
  (x => 256, y => 149),
  (x => 257, y => 149),
  (x => 258, y => 149),
  (x => 262, y => 149),
  (x => 263, y => 149),
  (x => 264, y => 149),
  (x => 265, y => 149),
  (x => 266, y => 149),
  (x => 267, y => 149),
  (x => 268, y => 149),
  (x => 269, y => 149),
  (x => 270, y => 149),
  (x => 271, y => 149),
  (x => 281, y => 149),
  (x => 282, y => 149),
  (x => 283, y => 149),
  (x => 284, y => 149),
  (x => 285, y => 149),
  (x => 286, y => 149),
  (x => 287, y => 149),
  (x => 288, y => 149),
  (x => 295, y => 149),
  (x => 296, y => 149),
  (x => 297, y => 149),
  (x => 298, y => 149),
  (x => 299, y => 149),
  (x => 300, y => 149),
  (x => 301, y => 149),
  (x => 323, y => 149),
  (x => 324, y => 149),
  (x => 325, y => 149),
  (x => 326, y => 149),
  (x => 327, y => 149),
  (x => 328, y => 149),
  (x => 329, y => 149),
  (x => 330, y => 149),
  (x => 351, y => 149),
  (x => 352, y => 149),
  (x => 353, y => 149),
  (x => 354, y => 149),
  (x => 355, y => 149),
  (x => 356, y => 149),
  (x => 357, y => 149),
  (x => 358, y => 149),
  (x => 364, y => 149),
  (x => 365, y => 149),
  (x => 366, y => 149),
  (x => 367, y => 149),
  (x => 368, y => 149),
  (x => 369, y => 149),
  (x => 370, y => 149),
  (x => 381, y => 149),
  (x => 382, y => 149),
  (x => 383, y => 149),
  (x => 384, y => 149),
  (x => 385, y => 149),
  (x => 386, y => 149),
  (x => 387, y => 149),
  (x => 396, y => 149),
  (x => 397, y => 149),
  (x => 398, y => 149),
  (x => 399, y => 149),
  (x => 400, y => 149),
  (x => 401, y => 149),
  (x => 402, y => 149),
  (x => 409, y => 149),
  (x => 410, y => 149),
  (x => 411, y => 149),
  (x => 412, y => 149),
  (x => 413, y => 149),
  (x => 414, y => 149),
  (x => 415, y => 149),
  (x => 424, y => 149),
  (x => 425, y => 149),
  (x => 426, y => 149),
  (x => 427, y => 149),
  (x => 428, y => 149),
  (x => 429, y => 149),
  (x => 430, y => 149),
  (x => 431, y => 149),
  (x => 432, y => 149),
  (x => 433, y => 149),
  (x => 434, y => 149),
  (x => 435, y => 149),
  (x => 436, y => 149),
  (x => 437, y => 149),
  (x => 438, y => 149),
  (x => 439, y => 149),
  (x => 162, y => 150),
  (x => 163, y => 150),
  (x => 164, y => 150),
  (x => 165, y => 150),
  (x => 166, y => 150),
  (x => 167, y => 150),
  (x => 168, y => 150),
  (x => 169, y => 150),
  (x => 179, y => 150),
  (x => 180, y => 150),
  (x => 181, y => 150),
  (x => 182, y => 150),
  (x => 183, y => 150),
  (x => 184, y => 150),
  (x => 185, y => 150),
  (x => 186, y => 150),
  (x => 187, y => 150),
  (x => 188, y => 150),
  (x => 189, y => 150),
  (x => 190, y => 150),
  (x => 191, y => 150),
  (x => 192, y => 150),
  (x => 193, y => 150),
  (x => 203, y => 150),
  (x => 216, y => 150),
  (x => 217, y => 150),
  (x => 218, y => 150),
  (x => 219, y => 150),
  (x => 220, y => 150),
  (x => 221, y => 150),
  (x => 231, y => 150),
  (x => 232, y => 150),
  (x => 233, y => 150),
  (x => 234, y => 150),
  (x => 235, y => 150),
  (x => 236, y => 150),
  (x => 237, y => 150),
  (x => 238, y => 150),
  (x => 239, y => 150),
  (x => 246, y => 150),
  (x => 247, y => 150),
  (x => 248, y => 150),
  (x => 249, y => 150),
  (x => 250, y => 150),
  (x => 251, y => 150),
  (x => 252, y => 150),
  (x => 253, y => 150),
  (x => 254, y => 150),
  (x => 255, y => 150),
  (x => 256, y => 150),
  (x => 257, y => 150),
  (x => 264, y => 150),
  (x => 265, y => 150),
  (x => 266, y => 150),
  (x => 267, y => 150),
  (x => 268, y => 150),
  (x => 269, y => 150),
  (x => 270, y => 150),
  (x => 271, y => 150),
  (x => 281, y => 150),
  (x => 282, y => 150),
  (x => 283, y => 150),
  (x => 284, y => 150),
  (x => 285, y => 150),
  (x => 286, y => 150),
  (x => 287, y => 150),
  (x => 296, y => 150),
  (x => 297, y => 150),
  (x => 298, y => 150),
  (x => 299, y => 150),
  (x => 300, y => 150),
  (x => 301, y => 150),
  (x => 323, y => 150),
  (x => 324, y => 150),
  (x => 325, y => 150),
  (x => 326, y => 150),
  (x => 327, y => 150),
  (x => 328, y => 150),
  (x => 329, y => 150),
  (x => 330, y => 150),
  (x => 351, y => 150),
  (x => 352, y => 150),
  (x => 353, y => 150),
  (x => 354, y => 150),
  (x => 355, y => 150),
  (x => 356, y => 150),
  (x => 357, y => 150),
  (x => 358, y => 150),
  (x => 365, y => 150),
  (x => 366, y => 150),
  (x => 367, y => 150),
  (x => 368, y => 150),
  (x => 369, y => 150),
  (x => 370, y => 150),
  (x => 381, y => 150),
  (x => 382, y => 150),
  (x => 383, y => 150),
  (x => 384, y => 150),
  (x => 385, y => 150),
  (x => 386, y => 150),
  (x => 387, y => 150),
  (x => 395, y => 150),
  (x => 396, y => 150),
  (x => 397, y => 150),
  (x => 398, y => 150),
  (x => 399, y => 150),
  (x => 400, y => 150),
  (x => 401, y => 150),
  (x => 410, y => 150),
  (x => 411, y => 150),
  (x => 412, y => 150),
  (x => 413, y => 150),
  (x => 414, y => 150),
  (x => 415, y => 150),
  (x => 416, y => 150),
  (x => 424, y => 150),
  (x => 425, y => 150),
  (x => 426, y => 150),
  (x => 427, y => 150),
  (x => 428, y => 150),
  (x => 429, y => 150),
  (x => 430, y => 150),
  (x => 431, y => 150),
  (x => 432, y => 150),
  (x => 433, y => 150),
  (x => 434, y => 150),
  (x => 435, y => 150),
  (x => 439, y => 150),
  (x => 162, y => 151),
  (x => 163, y => 151),
  (x => 164, y => 151),
  (x => 165, y => 151),
  (x => 166, y => 151),
  (x => 167, y => 151),
  (x => 168, y => 151),
  (x => 169, y => 151),
  (x => 179, y => 151),
  (x => 180, y => 151),
  (x => 181, y => 151),
  (x => 182, y => 151),
  (x => 183, y => 151),
  (x => 184, y => 151),
  (x => 185, y => 151),
  (x => 186, y => 151),
  (x => 187, y => 151),
  (x => 188, y => 151),
  (x => 189, y => 151),
  (x => 190, y => 151),
  (x => 191, y => 151),
  (x => 192, y => 151),
  (x => 193, y => 151),
  (x => 216, y => 151),
  (x => 217, y => 151),
  (x => 218, y => 151),
  (x => 219, y => 151),
  (x => 220, y => 151),
  (x => 221, y => 151),
  (x => 222, y => 151),
  (x => 231, y => 151),
  (x => 232, y => 151),
  (x => 233, y => 151),
  (x => 234, y => 151),
  (x => 235, y => 151),
  (x => 236, y => 151),
  (x => 237, y => 151),
  (x => 238, y => 151),
  (x => 239, y => 151),
  (x => 247, y => 151),
  (x => 248, y => 151),
  (x => 249, y => 151),
  (x => 250, y => 151),
  (x => 251, y => 151),
  (x => 252, y => 151),
  (x => 253, y => 151),
  (x => 254, y => 151),
  (x => 255, y => 151),
  (x => 256, y => 151),
  (x => 264, y => 151),
  (x => 265, y => 151),
  (x => 266, y => 151),
  (x => 267, y => 151),
  (x => 268, y => 151),
  (x => 269, y => 151),
  (x => 270, y => 151),
  (x => 271, y => 151),
  (x => 280, y => 151),
  (x => 281, y => 151),
  (x => 282, y => 151),
  (x => 283, y => 151),
  (x => 284, y => 151),
  (x => 285, y => 151),
  (x => 286, y => 151),
  (x => 296, y => 151),
  (x => 297, y => 151),
  (x => 298, y => 151),
  (x => 299, y => 151),
  (x => 300, y => 151),
  (x => 301, y => 151),
  (x => 323, y => 151),
  (x => 324, y => 151),
  (x => 325, y => 151),
  (x => 326, y => 151),
  (x => 327, y => 151),
  (x => 328, y => 151),
  (x => 329, y => 151),
  (x => 330, y => 151),
  (x => 351, y => 151),
  (x => 352, y => 151),
  (x => 353, y => 151),
  (x => 354, y => 151),
  (x => 355, y => 151),
  (x => 356, y => 151),
  (x => 357, y => 151),
  (x => 358, y => 151),
  (x => 365, y => 151),
  (x => 366, y => 151),
  (x => 367, y => 151),
  (x => 368, y => 151),
  (x => 369, y => 151),
  (x => 370, y => 151),
  (x => 371, y => 151),
  (x => 381, y => 151),
  (x => 382, y => 151),
  (x => 383, y => 151),
  (x => 384, y => 151),
  (x => 385, y => 151),
  (x => 386, y => 151),
  (x => 395, y => 151),
  (x => 396, y => 151),
  (x => 397, y => 151),
  (x => 398, y => 151),
  (x => 399, y => 151),
  (x => 400, y => 151),
  (x => 401, y => 151),
  (x => 411, y => 151),
  (x => 412, y => 151),
  (x => 413, y => 151),
  (x => 414, y => 151),
  (x => 415, y => 151),
  (x => 416, y => 151),
  (x => 424, y => 151),
  (x => 425, y => 151),
  (x => 426, y => 151),
  (x => 427, y => 151),
  (x => 428, y => 151),
  (x => 429, y => 151),
  (x => 430, y => 151),
  (x => 431, y => 151),
  (x => 432, y => 151),
  (x => 433, y => 151),
  (x => 162, y => 152),
  (x => 163, y => 152),
  (x => 164, y => 152),
  (x => 165, y => 152),
  (x => 166, y => 152),
  (x => 167, y => 152),
  (x => 168, y => 152),
  (x => 169, y => 152),
  (x => 179, y => 152),
  (x => 180, y => 152),
  (x => 181, y => 152),
  (x => 182, y => 152),
  (x => 183, y => 152),
  (x => 184, y => 152),
  (x => 185, y => 152),
  (x => 186, y => 152),
  (x => 187, y => 152),
  (x => 188, y => 152),
  (x => 189, y => 152),
  (x => 190, y => 152),
  (x => 191, y => 152),
  (x => 192, y => 152),
  (x => 193, y => 152),
  (x => 216, y => 152),
  (x => 217, y => 152),
  (x => 218, y => 152),
  (x => 219, y => 152),
  (x => 220, y => 152),
  (x => 221, y => 152),
  (x => 222, y => 152),
  (x => 231, y => 152),
  (x => 232, y => 152),
  (x => 233, y => 152),
  (x => 234, y => 152),
  (x => 235, y => 152),
  (x => 236, y => 152),
  (x => 237, y => 152),
  (x => 238, y => 152),
  (x => 248, y => 152),
  (x => 249, y => 152),
  (x => 250, y => 152),
  (x => 251, y => 152),
  (x => 252, y => 152),
  (x => 253, y => 152),
  (x => 254, y => 152),
  (x => 255, y => 152),
  (x => 265, y => 152),
  (x => 266, y => 152),
  (x => 267, y => 152),
  (x => 268, y => 152),
  (x => 269, y => 152),
  (x => 270, y => 152),
  (x => 271, y => 152),
  (x => 280, y => 152),
  (x => 281, y => 152),
  (x => 282, y => 152),
  (x => 283, y => 152),
  (x => 284, y => 152),
  (x => 285, y => 152),
  (x => 286, y => 152),
  (x => 297, y => 152),
  (x => 298, y => 152),
  (x => 299, y => 152),
  (x => 300, y => 152),
  (x => 301, y => 152),
  (x => 302, y => 152),
  (x => 323, y => 152),
  (x => 324, y => 152),
  (x => 325, y => 152),
  (x => 326, y => 152),
  (x => 327, y => 152),
  (x => 328, y => 152),
  (x => 329, y => 152),
  (x => 330, y => 152),
  (x => 351, y => 152),
  (x => 352, y => 152),
  (x => 353, y => 152),
  (x => 354, y => 152),
  (x => 355, y => 152),
  (x => 356, y => 152),
  (x => 357, y => 152),
  (x => 358, y => 152),
  (x => 365, y => 152),
  (x => 366, y => 152),
  (x => 367, y => 152),
  (x => 368, y => 152),
  (x => 369, y => 152),
  (x => 370, y => 152),
  (x => 371, y => 152),
  (x => 381, y => 152),
  (x => 382, y => 152),
  (x => 383, y => 152),
  (x => 384, y => 152),
  (x => 385, y => 152),
  (x => 386, y => 152),
  (x => 395, y => 152),
  (x => 396, y => 152),
  (x => 397, y => 152),
  (x => 398, y => 152),
  (x => 399, y => 152),
  (x => 400, y => 152),
  (x => 411, y => 152),
  (x => 412, y => 152),
  (x => 413, y => 152),
  (x => 414, y => 152),
  (x => 415, y => 152),
  (x => 416, y => 152),
  (x => 424, y => 152),
  (x => 425, y => 152),
  (x => 426, y => 152),
  (x => 427, y => 152),
  (x => 428, y => 152),
  (x => 429, y => 152),
  (x => 430, y => 152),
  (x => 431, y => 152),
  (x => 432, y => 152),
  (x => 162, y => 153),
  (x => 163, y => 153),
  (x => 164, y => 153),
  (x => 165, y => 153),
  (x => 166, y => 153),
  (x => 167, y => 153),
  (x => 168, y => 153),
  (x => 169, y => 153),
  (x => 179, y => 153),
  (x => 180, y => 153),
  (x => 181, y => 153),
  (x => 182, y => 153),
  (x => 183, y => 153),
  (x => 184, y => 153),
  (x => 185, y => 153),
  (x => 186, y => 153),
  (x => 187, y => 153),
  (x => 188, y => 153),
  (x => 189, y => 153),
  (x => 190, y => 153),
  (x => 191, y => 153),
  (x => 192, y => 153),
  (x => 193, y => 153),
  (x => 217, y => 153),
  (x => 218, y => 153),
  (x => 219, y => 153),
  (x => 220, y => 153),
  (x => 221, y => 153),
  (x => 222, y => 153),
  (x => 231, y => 153),
  (x => 232, y => 153),
  (x => 233, y => 153),
  (x => 234, y => 153),
  (x => 235, y => 153),
  (x => 236, y => 153),
  (x => 237, y => 153),
  (x => 238, y => 153),
  (x => 248, y => 153),
  (x => 249, y => 153),
  (x => 250, y => 153),
  (x => 251, y => 153),
  (x => 252, y => 153),
  (x => 253, y => 153),
  (x => 254, y => 153),
  (x => 255, y => 153),
  (x => 265, y => 153),
  (x => 266, y => 153),
  (x => 267, y => 153),
  (x => 268, y => 153),
  (x => 269, y => 153),
  (x => 270, y => 153),
  (x => 271, y => 153),
  (x => 280, y => 153),
  (x => 281, y => 153),
  (x => 282, y => 153),
  (x => 283, y => 153),
  (x => 284, y => 153),
  (x => 285, y => 153),
  (x => 297, y => 153),
  (x => 298, y => 153),
  (x => 299, y => 153),
  (x => 300, y => 153),
  (x => 301, y => 153),
  (x => 302, y => 153),
  (x => 323, y => 153),
  (x => 324, y => 153),
  (x => 325, y => 153),
  (x => 326, y => 153),
  (x => 327, y => 153),
  (x => 328, y => 153),
  (x => 329, y => 153),
  (x => 330, y => 153),
  (x => 351, y => 153),
  (x => 352, y => 153),
  (x => 353, y => 153),
  (x => 354, y => 153),
  (x => 355, y => 153),
  (x => 356, y => 153),
  (x => 357, y => 153),
  (x => 358, y => 153),
  (x => 365, y => 153),
  (x => 366, y => 153),
  (x => 367, y => 153),
  (x => 368, y => 153),
  (x => 369, y => 153),
  (x => 370, y => 153),
  (x => 371, y => 153),
  (x => 380, y => 153),
  (x => 381, y => 153),
  (x => 382, y => 153),
  (x => 383, y => 153),
  (x => 384, y => 153),
  (x => 385, y => 153),
  (x => 386, y => 153),
  (x => 394, y => 153),
  (x => 395, y => 153),
  (x => 396, y => 153),
  (x => 397, y => 153),
  (x => 398, y => 153),
  (x => 399, y => 153),
  (x => 400, y => 153),
  (x => 411, y => 153),
  (x => 412, y => 153),
  (x => 413, y => 153),
  (x => 414, y => 153),
  (x => 415, y => 153),
  (x => 416, y => 153),
  (x => 424, y => 153),
  (x => 425, y => 153),
  (x => 426, y => 153),
  (x => 427, y => 153),
  (x => 428, y => 153),
  (x => 429, y => 153),
  (x => 430, y => 153),
  (x => 431, y => 153),
  (x => 432, y => 153),
  (x => 162, y => 154),
  (x => 163, y => 154),
  (x => 164, y => 154),
  (x => 165, y => 154),
  (x => 166, y => 154),
  (x => 167, y => 154),
  (x => 168, y => 154),
  (x => 169, y => 154),
  (x => 179, y => 154),
  (x => 180, y => 154),
  (x => 181, y => 154),
  (x => 182, y => 154),
  (x => 183, y => 154),
  (x => 184, y => 154),
  (x => 185, y => 154),
  (x => 186, y => 154),
  (x => 187, y => 154),
  (x => 188, y => 154),
  (x => 189, y => 154),
  (x => 190, y => 154),
  (x => 191, y => 154),
  (x => 192, y => 154),
  (x => 193, y => 154),
  (x => 217, y => 154),
  (x => 218, y => 154),
  (x => 219, y => 154),
  (x => 220, y => 154),
  (x => 221, y => 154),
  (x => 222, y => 154),
  (x => 231, y => 154),
  (x => 232, y => 154),
  (x => 233, y => 154),
  (x => 234, y => 154),
  (x => 235, y => 154),
  (x => 236, y => 154),
  (x => 237, y => 154),
  (x => 248, y => 154),
  (x => 249, y => 154),
  (x => 250, y => 154),
  (x => 251, y => 154),
  (x => 252, y => 154),
  (x => 253, y => 154),
  (x => 254, y => 154),
  (x => 255, y => 154),
  (x => 265, y => 154),
  (x => 266, y => 154),
  (x => 267, y => 154),
  (x => 268, y => 154),
  (x => 269, y => 154),
  (x => 270, y => 154),
  (x => 271, y => 154),
  (x => 280, y => 154),
  (x => 281, y => 154),
  (x => 282, y => 154),
  (x => 283, y => 154),
  (x => 284, y => 154),
  (x => 285, y => 154),
  (x => 297, y => 154),
  (x => 298, y => 154),
  (x => 299, y => 154),
  (x => 300, y => 154),
  (x => 301, y => 154),
  (x => 302, y => 154),
  (x => 323, y => 154),
  (x => 324, y => 154),
  (x => 325, y => 154),
  (x => 326, y => 154),
  (x => 327, y => 154),
  (x => 328, y => 154),
  (x => 329, y => 154),
  (x => 330, y => 154),
  (x => 351, y => 154),
  (x => 352, y => 154),
  (x => 353, y => 154),
  (x => 354, y => 154),
  (x => 355, y => 154),
  (x => 356, y => 154),
  (x => 357, y => 154),
  (x => 358, y => 154),
  (x => 366, y => 154),
  (x => 367, y => 154),
  (x => 368, y => 154),
  (x => 369, y => 154),
  (x => 370, y => 154),
  (x => 371, y => 154),
  (x => 380, y => 154),
  (x => 381, y => 154),
  (x => 382, y => 154),
  (x => 383, y => 154),
  (x => 384, y => 154),
  (x => 385, y => 154),
  (x => 386, y => 154),
  (x => 394, y => 154),
  (x => 395, y => 154),
  (x => 396, y => 154),
  (x => 397, y => 154),
  (x => 398, y => 154),
  (x => 399, y => 154),
  (x => 400, y => 154),
  (x => 411, y => 154),
  (x => 412, y => 154),
  (x => 413, y => 154),
  (x => 414, y => 154),
  (x => 415, y => 154),
  (x => 416, y => 154),
  (x => 417, y => 154),
  (x => 424, y => 154),
  (x => 425, y => 154),
  (x => 426, y => 154),
  (x => 427, y => 154),
  (x => 428, y => 154),
  (x => 429, y => 154),
  (x => 430, y => 154),
  (x => 431, y => 154),
  (x => 162, y => 155),
  (x => 163, y => 155),
  (x => 164, y => 155),
  (x => 165, y => 155),
  (x => 166, y => 155),
  (x => 167, y => 155),
  (x => 168, y => 155),
  (x => 169, y => 155),
  (x => 179, y => 155),
  (x => 180, y => 155),
  (x => 181, y => 155),
  (x => 182, y => 155),
  (x => 183, y => 155),
  (x => 184, y => 155),
  (x => 185, y => 155),
  (x => 186, y => 155),
  (x => 187, y => 155),
  (x => 188, y => 155),
  (x => 189, y => 155),
  (x => 190, y => 155),
  (x => 191, y => 155),
  (x => 192, y => 155),
  (x => 193, y => 155),
  (x => 216, y => 155),
  (x => 217, y => 155),
  (x => 218, y => 155),
  (x => 219, y => 155),
  (x => 220, y => 155),
  (x => 221, y => 155),
  (x => 222, y => 155),
  (x => 231, y => 155),
  (x => 232, y => 155),
  (x => 233, y => 155),
  (x => 234, y => 155),
  (x => 235, y => 155),
  (x => 236, y => 155),
  (x => 237, y => 155),
  (x => 248, y => 155),
  (x => 249, y => 155),
  (x => 250, y => 155),
  (x => 251, y => 155),
  (x => 252, y => 155),
  (x => 253, y => 155),
  (x => 254, y => 155),
  (x => 266, y => 155),
  (x => 267, y => 155),
  (x => 268, y => 155),
  (x => 269, y => 155),
  (x => 270, y => 155),
  (x => 271, y => 155),
  (x => 272, y => 155),
  (x => 279, y => 155),
  (x => 280, y => 155),
  (x => 281, y => 155),
  (x => 282, y => 155),
  (x => 283, y => 155),
  (x => 284, y => 155),
  (x => 285, y => 155),
  (x => 297, y => 155),
  (x => 298, y => 155),
  (x => 299, y => 155),
  (x => 300, y => 155),
  (x => 301, y => 155),
  (x => 302, y => 155),
  (x => 323, y => 155),
  (x => 324, y => 155),
  (x => 325, y => 155),
  (x => 326, y => 155),
  (x => 327, y => 155),
  (x => 328, y => 155),
  (x => 329, y => 155),
  (x => 330, y => 155),
  (x => 351, y => 155),
  (x => 352, y => 155),
  (x => 353, y => 155),
  (x => 354, y => 155),
  (x => 355, y => 155),
  (x => 356, y => 155),
  (x => 357, y => 155),
  (x => 358, y => 155),
  (x => 366, y => 155),
  (x => 367, y => 155),
  (x => 368, y => 155),
  (x => 369, y => 155),
  (x => 370, y => 155),
  (x => 371, y => 155),
  (x => 372, y => 155),
  (x => 380, y => 155),
  (x => 381, y => 155),
  (x => 382, y => 155),
  (x => 383, y => 155),
  (x => 384, y => 155),
  (x => 385, y => 155),
  (x => 394, y => 155),
  (x => 395, y => 155),
  (x => 396, y => 155),
  (x => 397, y => 155),
  (x => 398, y => 155),
  (x => 399, y => 155),
  (x => 412, y => 155),
  (x => 413, y => 155),
  (x => 414, y => 155),
  (x => 415, y => 155),
  (x => 416, y => 155),
  (x => 417, y => 155),
  (x => 424, y => 155),
  (x => 425, y => 155),
  (x => 426, y => 155),
  (x => 427, y => 155),
  (x => 428, y => 155),
  (x => 429, y => 155),
  (x => 430, y => 155),
  (x => 431, y => 155),
  (x => 162, y => 156),
  (x => 163, y => 156),
  (x => 164, y => 156),
  (x => 165, y => 156),
  (x => 166, y => 156),
  (x => 167, y => 156),
  (x => 168, y => 156),
  (x => 169, y => 156),
  (x => 179, y => 156),
  (x => 180, y => 156),
  (x => 181, y => 156),
  (x => 182, y => 156),
  (x => 183, y => 156),
  (x => 184, y => 156),
  (x => 185, y => 156),
  (x => 186, y => 156),
  (x => 187, y => 156),
  (x => 188, y => 156),
  (x => 189, y => 156),
  (x => 190, y => 156),
  (x => 191, y => 156),
  (x => 192, y => 156),
  (x => 193, y => 156),
  (x => 212, y => 156),
  (x => 213, y => 156),
  (x => 214, y => 156),
  (x => 215, y => 156),
  (x => 216, y => 156),
  (x => 217, y => 156),
  (x => 218, y => 156),
  (x => 219, y => 156),
  (x => 220, y => 156),
  (x => 221, y => 156),
  (x => 222, y => 156),
  (x => 231, y => 156),
  (x => 232, y => 156),
  (x => 233, y => 156),
  (x => 234, y => 156),
  (x => 235, y => 156),
  (x => 236, y => 156),
  (x => 237, y => 156),
  (x => 248, y => 156),
  (x => 249, y => 156),
  (x => 250, y => 156),
  (x => 251, y => 156),
  (x => 252, y => 156),
  (x => 253, y => 156),
  (x => 254, y => 156),
  (x => 266, y => 156),
  (x => 267, y => 156),
  (x => 268, y => 156),
  (x => 269, y => 156),
  (x => 270, y => 156),
  (x => 271, y => 156),
  (x => 272, y => 156),
  (x => 279, y => 156),
  (x => 280, y => 156),
  (x => 281, y => 156),
  (x => 282, y => 156),
  (x => 283, y => 156),
  (x => 284, y => 156),
  (x => 285, y => 156),
  (x => 297, y => 156),
  (x => 298, y => 156),
  (x => 299, y => 156),
  (x => 300, y => 156),
  (x => 301, y => 156),
  (x => 302, y => 156),
  (x => 323, y => 156),
  (x => 324, y => 156),
  (x => 325, y => 156),
  (x => 326, y => 156),
  (x => 327, y => 156),
  (x => 328, y => 156),
  (x => 329, y => 156),
  (x => 330, y => 156),
  (x => 351, y => 156),
  (x => 352, y => 156),
  (x => 353, y => 156),
  (x => 354, y => 156),
  (x => 355, y => 156),
  (x => 356, y => 156),
  (x => 357, y => 156),
  (x => 358, y => 156),
  (x => 366, y => 156),
  (x => 367, y => 156),
  (x => 368, y => 156),
  (x => 369, y => 156),
  (x => 370, y => 156),
  (x => 371, y => 156),
  (x => 372, y => 156),
  (x => 380, y => 156),
  (x => 381, y => 156),
  (x => 382, y => 156),
  (x => 383, y => 156),
  (x => 384, y => 156),
  (x => 385, y => 156),
  (x => 394, y => 156),
  (x => 395, y => 156),
  (x => 396, y => 156),
  (x => 397, y => 156),
  (x => 398, y => 156),
  (x => 399, y => 156),
  (x => 412, y => 156),
  (x => 413, y => 156),
  (x => 414, y => 156),
  (x => 415, y => 156),
  (x => 416, y => 156),
  (x => 417, y => 156),
  (x => 424, y => 156),
  (x => 425, y => 156),
  (x => 426, y => 156),
  (x => 427, y => 156),
  (x => 428, y => 156),
  (x => 429, y => 156),
  (x => 430, y => 156),
  (x => 431, y => 156),
  (x => 162, y => 157),
  (x => 163, y => 157),
  (x => 164, y => 157),
  (x => 165, y => 157),
  (x => 166, y => 157),
  (x => 167, y => 157),
  (x => 168, y => 157),
  (x => 169, y => 157),
  (x => 179, y => 157),
  (x => 180, y => 157),
  (x => 181, y => 157),
  (x => 182, y => 157),
  (x => 183, y => 157),
  (x => 184, y => 157),
  (x => 185, y => 157),
  (x => 186, y => 157),
  (x => 187, y => 157),
  (x => 188, y => 157),
  (x => 189, y => 157),
  (x => 190, y => 157),
  (x => 191, y => 157),
  (x => 192, y => 157),
  (x => 193, y => 157),
  (x => 207, y => 157),
  (x => 208, y => 157),
  (x => 209, y => 157),
  (x => 210, y => 157),
  (x => 211, y => 157),
  (x => 212, y => 157),
  (x => 213, y => 157),
  (x => 214, y => 157),
  (x => 215, y => 157),
  (x => 216, y => 157),
  (x => 217, y => 157),
  (x => 218, y => 157),
  (x => 219, y => 157),
  (x => 220, y => 157),
  (x => 221, y => 157),
  (x => 222, y => 157),
  (x => 231, y => 157),
  (x => 232, y => 157),
  (x => 233, y => 157),
  (x => 234, y => 157),
  (x => 235, y => 157),
  (x => 236, y => 157),
  (x => 237, y => 157),
  (x => 248, y => 157),
  (x => 249, y => 157),
  (x => 250, y => 157),
  (x => 251, y => 157),
  (x => 252, y => 157),
  (x => 253, y => 157),
  (x => 254, y => 157),
  (x => 266, y => 157),
  (x => 267, y => 157),
  (x => 268, y => 157),
  (x => 269, y => 157),
  (x => 270, y => 157),
  (x => 271, y => 157),
  (x => 272, y => 157),
  (x => 279, y => 157),
  (x => 280, y => 157),
  (x => 281, y => 157),
  (x => 282, y => 157),
  (x => 283, y => 157),
  (x => 284, y => 157),
  (x => 285, y => 157),
  (x => 297, y => 157),
  (x => 298, y => 157),
  (x => 299, y => 157),
  (x => 300, y => 157),
  (x => 301, y => 157),
  (x => 302, y => 157),
  (x => 323, y => 157),
  (x => 324, y => 157),
  (x => 325, y => 157),
  (x => 326, y => 157),
  (x => 327, y => 157),
  (x => 328, y => 157),
  (x => 329, y => 157),
  (x => 330, y => 157),
  (x => 351, y => 157),
  (x => 352, y => 157),
  (x => 353, y => 157),
  (x => 354, y => 157),
  (x => 355, y => 157),
  (x => 356, y => 157),
  (x => 357, y => 157),
  (x => 358, y => 157),
  (x => 366, y => 157),
  (x => 367, y => 157),
  (x => 368, y => 157),
  (x => 369, y => 157),
  (x => 370, y => 157),
  (x => 371, y => 157),
  (x => 372, y => 157),
  (x => 380, y => 157),
  (x => 381, y => 157),
  (x => 382, y => 157),
  (x => 383, y => 157),
  (x => 384, y => 157),
  (x => 385, y => 157),
  (x => 394, y => 157),
  (x => 395, y => 157),
  (x => 396, y => 157),
  (x => 397, y => 157),
  (x => 398, y => 157),
  (x => 399, y => 157),
  (x => 412, y => 157),
  (x => 413, y => 157),
  (x => 414, y => 157),
  (x => 415, y => 157),
  (x => 416, y => 157),
  (x => 417, y => 157),
  (x => 424, y => 157),
  (x => 425, y => 157),
  (x => 426, y => 157),
  (x => 427, y => 157),
  (x => 428, y => 157),
  (x => 429, y => 157),
  (x => 430, y => 157),
  (x => 162, y => 158),
  (x => 163, y => 158),
  (x => 164, y => 158),
  (x => 165, y => 158),
  (x => 166, y => 158),
  (x => 167, y => 158),
  (x => 168, y => 158),
  (x => 169, y => 158),
  (x => 187, y => 158),
  (x => 188, y => 158),
  (x => 189, y => 158),
  (x => 190, y => 158),
  (x => 191, y => 158),
  (x => 192, y => 158),
  (x => 193, y => 158),
  (x => 205, y => 158),
  (x => 206, y => 158),
  (x => 207, y => 158),
  (x => 208, y => 158),
  (x => 209, y => 158),
  (x => 210, y => 158),
  (x => 211, y => 158),
  (x => 212, y => 158),
  (x => 213, y => 158),
  (x => 214, y => 158),
  (x => 215, y => 158),
  (x => 216, y => 158),
  (x => 217, y => 158),
  (x => 218, y => 158),
  (x => 219, y => 158),
  (x => 220, y => 158),
  (x => 221, y => 158),
  (x => 222, y => 158),
  (x => 231, y => 158),
  (x => 232, y => 158),
  (x => 233, y => 158),
  (x => 234, y => 158),
  (x => 235, y => 158),
  (x => 236, y => 158),
  (x => 237, y => 158),
  (x => 248, y => 158),
  (x => 249, y => 158),
  (x => 250, y => 158),
  (x => 251, y => 158),
  (x => 252, y => 158),
  (x => 253, y => 158),
  (x => 254, y => 158),
  (x => 266, y => 158),
  (x => 267, y => 158),
  (x => 268, y => 158),
  (x => 269, y => 158),
  (x => 270, y => 158),
  (x => 271, y => 158),
  (x => 272, y => 158),
  (x => 279, y => 158),
  (x => 280, y => 158),
  (x => 281, y => 158),
  (x => 282, y => 158),
  (x => 283, y => 158),
  (x => 284, y => 158),
  (x => 285, y => 158),
  (x => 286, y => 158),
  (x => 287, y => 158),
  (x => 288, y => 158),
  (x => 289, y => 158),
  (x => 290, y => 158),
  (x => 291, y => 158),
  (x => 292, y => 158),
  (x => 293, y => 158),
  (x => 294, y => 158),
  (x => 295, y => 158),
  (x => 296, y => 158),
  (x => 297, y => 158),
  (x => 298, y => 158),
  (x => 299, y => 158),
  (x => 300, y => 158),
  (x => 301, y => 158),
  (x => 302, y => 158),
  (x => 323, y => 158),
  (x => 324, y => 158),
  (x => 325, y => 158),
  (x => 326, y => 158),
  (x => 327, y => 158),
  (x => 328, y => 158),
  (x => 329, y => 158),
  (x => 330, y => 158),
  (x => 351, y => 158),
  (x => 352, y => 158),
  (x => 353, y => 158),
  (x => 354, y => 158),
  (x => 355, y => 158),
  (x => 356, y => 158),
  (x => 357, y => 158),
  (x => 358, y => 158),
  (x => 367, y => 158),
  (x => 368, y => 158),
  (x => 369, y => 158),
  (x => 370, y => 158),
  (x => 371, y => 158),
  (x => 372, y => 158),
  (x => 379, y => 158),
  (x => 380, y => 158),
  (x => 381, y => 158),
  (x => 382, y => 158),
  (x => 383, y => 158),
  (x => 384, y => 158),
  (x => 385, y => 158),
  (x => 394, y => 158),
  (x => 395, y => 158),
  (x => 396, y => 158),
  (x => 397, y => 158),
  (x => 398, y => 158),
  (x => 399, y => 158),
  (x => 400, y => 158),
  (x => 401, y => 158),
  (x => 402, y => 158),
  (x => 403, y => 158),
  (x => 404, y => 158),
  (x => 405, y => 158),
  (x => 406, y => 158),
  (x => 407, y => 158),
  (x => 408, y => 158),
  (x => 409, y => 158),
  (x => 410, y => 158),
  (x => 411, y => 158),
  (x => 412, y => 158),
  (x => 413, y => 158),
  (x => 414, y => 158),
  (x => 415, y => 158),
  (x => 416, y => 158),
  (x => 417, y => 158),
  (x => 424, y => 158),
  (x => 425, y => 158),
  (x => 426, y => 158),
  (x => 427, y => 158),
  (x => 428, y => 158),
  (x => 429, y => 158),
  (x => 430, y => 158),
  (x => 162, y => 159),
  (x => 163, y => 159),
  (x => 164, y => 159),
  (x => 165, y => 159),
  (x => 166, y => 159),
  (x => 167, y => 159),
  (x => 168, y => 159),
  (x => 169, y => 159),
  (x => 187, y => 159),
  (x => 188, y => 159),
  (x => 189, y => 159),
  (x => 190, y => 159),
  (x => 191, y => 159),
  (x => 192, y => 159),
  (x => 193, y => 159),
  (x => 203, y => 159),
  (x => 204, y => 159),
  (x => 205, y => 159),
  (x => 206, y => 159),
  (x => 207, y => 159),
  (x => 208, y => 159),
  (x => 209, y => 159),
  (x => 210, y => 159),
  (x => 211, y => 159),
  (x => 212, y => 159),
  (x => 213, y => 159),
  (x => 214, y => 159),
  (x => 215, y => 159),
  (x => 216, y => 159),
  (x => 217, y => 159),
  (x => 218, y => 159),
  (x => 219, y => 159),
  (x => 220, y => 159),
  (x => 221, y => 159),
  (x => 222, y => 159),
  (x => 231, y => 159),
  (x => 232, y => 159),
  (x => 233, y => 159),
  (x => 234, y => 159),
  (x => 235, y => 159),
  (x => 236, y => 159),
  (x => 237, y => 159),
  (x => 248, y => 159),
  (x => 249, y => 159),
  (x => 250, y => 159),
  (x => 251, y => 159),
  (x => 252, y => 159),
  (x => 253, y => 159),
  (x => 254, y => 159),
  (x => 266, y => 159),
  (x => 267, y => 159),
  (x => 268, y => 159),
  (x => 269, y => 159),
  (x => 270, y => 159),
  (x => 271, y => 159),
  (x => 272, y => 159),
  (x => 279, y => 159),
  (x => 280, y => 159),
  (x => 281, y => 159),
  (x => 282, y => 159),
  (x => 283, y => 159),
  (x => 284, y => 159),
  (x => 285, y => 159),
  (x => 286, y => 159),
  (x => 287, y => 159),
  (x => 288, y => 159),
  (x => 289, y => 159),
  (x => 290, y => 159),
  (x => 291, y => 159),
  (x => 292, y => 159),
  (x => 293, y => 159),
  (x => 294, y => 159),
  (x => 295, y => 159),
  (x => 296, y => 159),
  (x => 297, y => 159),
  (x => 298, y => 159),
  (x => 299, y => 159),
  (x => 300, y => 159),
  (x => 301, y => 159),
  (x => 302, y => 159),
  (x => 324, y => 159),
  (x => 325, y => 159),
  (x => 326, y => 159),
  (x => 327, y => 159),
  (x => 328, y => 159),
  (x => 329, y => 159),
  (x => 330, y => 159),
  (x => 351, y => 159),
  (x => 352, y => 159),
  (x => 353, y => 159),
  (x => 354, y => 159),
  (x => 355, y => 159),
  (x => 356, y => 159),
  (x => 357, y => 159),
  (x => 367, y => 159),
  (x => 368, y => 159),
  (x => 369, y => 159),
  (x => 370, y => 159),
  (x => 371, y => 159),
  (x => 372, y => 159),
  (x => 379, y => 159),
  (x => 380, y => 159),
  (x => 381, y => 159),
  (x => 382, y => 159),
  (x => 383, y => 159),
  (x => 384, y => 159),
  (x => 393, y => 159),
  (x => 394, y => 159),
  (x => 395, y => 159),
  (x => 396, y => 159),
  (x => 397, y => 159),
  (x => 398, y => 159),
  (x => 399, y => 159),
  (x => 400, y => 159),
  (x => 401, y => 159),
  (x => 402, y => 159),
  (x => 403, y => 159),
  (x => 404, y => 159),
  (x => 405, y => 159),
  (x => 406, y => 159),
  (x => 407, y => 159),
  (x => 408, y => 159),
  (x => 409, y => 159),
  (x => 410, y => 159),
  (x => 411, y => 159),
  (x => 412, y => 159),
  (x => 413, y => 159),
  (x => 414, y => 159),
  (x => 415, y => 159),
  (x => 416, y => 159),
  (x => 417, y => 159),
  (x => 424, y => 159),
  (x => 425, y => 159),
  (x => 426, y => 159),
  (x => 427, y => 159),
  (x => 428, y => 159),
  (x => 429, y => 159),
  (x => 430, y => 159),
  (x => 163, y => 160),
  (x => 164, y => 160),
  (x => 165, y => 160),
  (x => 166, y => 160),
  (x => 167, y => 160),
  (x => 168, y => 160),
  (x => 169, y => 160),
  (x => 187, y => 160),
  (x => 188, y => 160),
  (x => 189, y => 160),
  (x => 190, y => 160),
  (x => 191, y => 160),
  (x => 192, y => 160),
  (x => 193, y => 160),
  (x => 202, y => 160),
  (x => 203, y => 160),
  (x => 204, y => 160),
  (x => 205, y => 160),
  (x => 206, y => 160),
  (x => 207, y => 160),
  (x => 208, y => 160),
  (x => 209, y => 160),
  (x => 210, y => 160),
  (x => 211, y => 160),
  (x => 212, y => 160),
  (x => 213, y => 160),
  (x => 214, y => 160),
  (x => 215, y => 160),
  (x => 216, y => 160),
  (x => 217, y => 160),
  (x => 218, y => 160),
  (x => 219, y => 160),
  (x => 220, y => 160),
  (x => 221, y => 160),
  (x => 222, y => 160),
  (x => 231, y => 160),
  (x => 232, y => 160),
  (x => 233, y => 160),
  (x => 234, y => 160),
  (x => 235, y => 160),
  (x => 236, y => 160),
  (x => 237, y => 160),
  (x => 248, y => 160),
  (x => 249, y => 160),
  (x => 250, y => 160),
  (x => 251, y => 160),
  (x => 252, y => 160),
  (x => 253, y => 160),
  (x => 254, y => 160),
  (x => 266, y => 160),
  (x => 267, y => 160),
  (x => 268, y => 160),
  (x => 269, y => 160),
  (x => 270, y => 160),
  (x => 271, y => 160),
  (x => 272, y => 160),
  (x => 279, y => 160),
  (x => 280, y => 160),
  (x => 281, y => 160),
  (x => 282, y => 160),
  (x => 283, y => 160),
  (x => 284, y => 160),
  (x => 285, y => 160),
  (x => 286, y => 160),
  (x => 287, y => 160),
  (x => 288, y => 160),
  (x => 289, y => 160),
  (x => 290, y => 160),
  (x => 291, y => 160),
  (x => 292, y => 160),
  (x => 293, y => 160),
  (x => 294, y => 160),
  (x => 295, y => 160),
  (x => 296, y => 160),
  (x => 297, y => 160),
  (x => 298, y => 160),
  (x => 299, y => 160),
  (x => 300, y => 160),
  (x => 301, y => 160),
  (x => 302, y => 160),
  (x => 324, y => 160),
  (x => 325, y => 160),
  (x => 326, y => 160),
  (x => 327, y => 160),
  (x => 328, y => 160),
  (x => 329, y => 160),
  (x => 330, y => 160),
  (x => 331, y => 160),
  (x => 351, y => 160),
  (x => 352, y => 160),
  (x => 353, y => 160),
  (x => 354, y => 160),
  (x => 355, y => 160),
  (x => 356, y => 160),
  (x => 357, y => 160),
  (x => 367, y => 160),
  (x => 368, y => 160),
  (x => 369, y => 160),
  (x => 370, y => 160),
  (x => 371, y => 160),
  (x => 372, y => 160),
  (x => 373, y => 160),
  (x => 379, y => 160),
  (x => 380, y => 160),
  (x => 381, y => 160),
  (x => 382, y => 160),
  (x => 383, y => 160),
  (x => 384, y => 160),
  (x => 393, y => 160),
  (x => 394, y => 160),
  (x => 395, y => 160),
  (x => 396, y => 160),
  (x => 397, y => 160),
  (x => 398, y => 160),
  (x => 399, y => 160),
  (x => 400, y => 160),
  (x => 401, y => 160),
  (x => 402, y => 160),
  (x => 403, y => 160),
  (x => 404, y => 160),
  (x => 405, y => 160),
  (x => 406, y => 160),
  (x => 407, y => 160),
  (x => 408, y => 160),
  (x => 409, y => 160),
  (x => 410, y => 160),
  (x => 411, y => 160),
  (x => 412, y => 160),
  (x => 413, y => 160),
  (x => 414, y => 160),
  (x => 415, y => 160),
  (x => 416, y => 160),
  (x => 417, y => 160),
  (x => 424, y => 160),
  (x => 425, y => 160),
  (x => 426, y => 160),
  (x => 427, y => 160),
  (x => 428, y => 160),
  (x => 429, y => 160),
  (x => 430, y => 160),
  (x => 163, y => 161),
  (x => 164, y => 161),
  (x => 165, y => 161),
  (x => 166, y => 161),
  (x => 167, y => 161),
  (x => 168, y => 161),
  (x => 169, y => 161),
  (x => 170, y => 161),
  (x => 187, y => 161),
  (x => 188, y => 161),
  (x => 189, y => 161),
  (x => 190, y => 161),
  (x => 191, y => 161),
  (x => 192, y => 161),
  (x => 193, y => 161),
  (x => 202, y => 161),
  (x => 203, y => 161),
  (x => 204, y => 161),
  (x => 205, y => 161),
  (x => 206, y => 161),
  (x => 207, y => 161),
  (x => 208, y => 161),
  (x => 209, y => 161),
  (x => 210, y => 161),
  (x => 217, y => 161),
  (x => 218, y => 161),
  (x => 219, y => 161),
  (x => 220, y => 161),
  (x => 221, y => 161),
  (x => 222, y => 161),
  (x => 231, y => 161),
  (x => 232, y => 161),
  (x => 233, y => 161),
  (x => 234, y => 161),
  (x => 235, y => 161),
  (x => 236, y => 161),
  (x => 237, y => 161),
  (x => 248, y => 161),
  (x => 249, y => 161),
  (x => 250, y => 161),
  (x => 251, y => 161),
  (x => 252, y => 161),
  (x => 253, y => 161),
  (x => 254, y => 161),
  (x => 266, y => 161),
  (x => 267, y => 161),
  (x => 268, y => 161),
  (x => 269, y => 161),
  (x => 270, y => 161),
  (x => 271, y => 161),
  (x => 272, y => 161),
  (x => 279, y => 161),
  (x => 280, y => 161),
  (x => 281, y => 161),
  (x => 282, y => 161),
  (x => 283, y => 161),
  (x => 284, y => 161),
  (x => 285, y => 161),
  (x => 286, y => 161),
  (x => 287, y => 161),
  (x => 288, y => 161),
  (x => 289, y => 161),
  (x => 290, y => 161),
  (x => 291, y => 161),
  (x => 292, y => 161),
  (x => 293, y => 161),
  (x => 294, y => 161),
  (x => 295, y => 161),
  (x => 296, y => 161),
  (x => 297, y => 161),
  (x => 298, y => 161),
  (x => 299, y => 161),
  (x => 300, y => 161),
  (x => 301, y => 161),
  (x => 302, y => 161),
  (x => 324, y => 161),
  (x => 325, y => 161),
  (x => 326, y => 161),
  (x => 327, y => 161),
  (x => 328, y => 161),
  (x => 329, y => 161),
  (x => 330, y => 161),
  (x => 331, y => 161),
  (x => 350, y => 161),
  (x => 351, y => 161),
  (x => 352, y => 161),
  (x => 353, y => 161),
  (x => 354, y => 161),
  (x => 355, y => 161),
  (x => 356, y => 161),
  (x => 357, y => 161),
  (x => 367, y => 161),
  (x => 368, y => 161),
  (x => 369, y => 161),
  (x => 370, y => 161),
  (x => 371, y => 161),
  (x => 372, y => 161),
  (x => 373, y => 161),
  (x => 379, y => 161),
  (x => 380, y => 161),
  (x => 381, y => 161),
  (x => 382, y => 161),
  (x => 383, y => 161),
  (x => 384, y => 161),
  (x => 393, y => 161),
  (x => 394, y => 161),
  (x => 395, y => 161),
  (x => 396, y => 161),
  (x => 397, y => 161),
  (x => 398, y => 161),
  (x => 399, y => 161),
  (x => 400, y => 161),
  (x => 401, y => 161),
  (x => 402, y => 161),
  (x => 403, y => 161),
  (x => 404, y => 161),
  (x => 405, y => 161),
  (x => 406, y => 161),
  (x => 407, y => 161),
  (x => 408, y => 161),
  (x => 409, y => 161),
  (x => 410, y => 161),
  (x => 411, y => 161),
  (x => 412, y => 161),
  (x => 413, y => 161),
  (x => 414, y => 161),
  (x => 415, y => 161),
  (x => 416, y => 161),
  (x => 417, y => 161),
  (x => 424, y => 161),
  (x => 425, y => 161),
  (x => 426, y => 161),
  (x => 427, y => 161),
  (x => 428, y => 161),
  (x => 429, y => 161),
  (x => 430, y => 161),
  (x => 163, y => 162),
  (x => 164, y => 162),
  (x => 165, y => 162),
  (x => 166, y => 162),
  (x => 167, y => 162),
  (x => 168, y => 162),
  (x => 169, y => 162),
  (x => 170, y => 162),
  (x => 187, y => 162),
  (x => 188, y => 162),
  (x => 189, y => 162),
  (x => 190, y => 162),
  (x => 191, y => 162),
  (x => 192, y => 162),
  (x => 193, y => 162),
  (x => 201, y => 162),
  (x => 202, y => 162),
  (x => 203, y => 162),
  (x => 204, y => 162),
  (x => 205, y => 162),
  (x => 206, y => 162),
  (x => 207, y => 162),
  (x => 208, y => 162),
  (x => 217, y => 162),
  (x => 218, y => 162),
  (x => 219, y => 162),
  (x => 220, y => 162),
  (x => 221, y => 162),
  (x => 222, y => 162),
  (x => 231, y => 162),
  (x => 232, y => 162),
  (x => 233, y => 162),
  (x => 234, y => 162),
  (x => 235, y => 162),
  (x => 236, y => 162),
  (x => 237, y => 162),
  (x => 248, y => 162),
  (x => 249, y => 162),
  (x => 250, y => 162),
  (x => 251, y => 162),
  (x => 252, y => 162),
  (x => 253, y => 162),
  (x => 254, y => 162),
  (x => 266, y => 162),
  (x => 267, y => 162),
  (x => 268, y => 162),
  (x => 269, y => 162),
  (x => 270, y => 162),
  (x => 271, y => 162),
  (x => 272, y => 162),
  (x => 279, y => 162),
  (x => 280, y => 162),
  (x => 281, y => 162),
  (x => 282, y => 162),
  (x => 283, y => 162),
  (x => 284, y => 162),
  (x => 285, y => 162),
  (x => 286, y => 162),
  (x => 287, y => 162),
  (x => 288, y => 162),
  (x => 289, y => 162),
  (x => 290, y => 162),
  (x => 291, y => 162),
  (x => 292, y => 162),
  (x => 293, y => 162),
  (x => 294, y => 162),
  (x => 295, y => 162),
  (x => 296, y => 162),
  (x => 297, y => 162),
  (x => 298, y => 162),
  (x => 299, y => 162),
  (x => 300, y => 162),
  (x => 301, y => 162),
  (x => 302, y => 162),
  (x => 324, y => 162),
  (x => 325, y => 162),
  (x => 326, y => 162),
  (x => 327, y => 162),
  (x => 328, y => 162),
  (x => 329, y => 162),
  (x => 330, y => 162),
  (x => 331, y => 162),
  (x => 350, y => 162),
  (x => 351, y => 162),
  (x => 352, y => 162),
  (x => 353, y => 162),
  (x => 354, y => 162),
  (x => 355, y => 162),
  (x => 356, y => 162),
  (x => 357, y => 162),
  (x => 368, y => 162),
  (x => 369, y => 162),
  (x => 370, y => 162),
  (x => 371, y => 162),
  (x => 372, y => 162),
  (x => 373, y => 162),
  (x => 378, y => 162),
  (x => 379, y => 162),
  (x => 380, y => 162),
  (x => 381, y => 162),
  (x => 382, y => 162),
  (x => 383, y => 162),
  (x => 393, y => 162),
  (x => 394, y => 162),
  (x => 395, y => 162),
  (x => 396, y => 162),
  (x => 397, y => 162),
  (x => 398, y => 162),
  (x => 399, y => 162),
  (x => 400, y => 162),
  (x => 401, y => 162),
  (x => 402, y => 162),
  (x => 403, y => 162),
  (x => 404, y => 162),
  (x => 405, y => 162),
  (x => 406, y => 162),
  (x => 407, y => 162),
  (x => 408, y => 162),
  (x => 409, y => 162),
  (x => 410, y => 162),
  (x => 411, y => 162),
  (x => 412, y => 162),
  (x => 413, y => 162),
  (x => 414, y => 162),
  (x => 415, y => 162),
  (x => 416, y => 162),
  (x => 417, y => 162),
  (x => 424, y => 162),
  (x => 425, y => 162),
  (x => 426, y => 162),
  (x => 427, y => 162),
  (x => 428, y => 162),
  (x => 429, y => 162),
  (x => 430, y => 162),
  (x => 163, y => 163),
  (x => 164, y => 163),
  (x => 165, y => 163),
  (x => 166, y => 163),
  (x => 167, y => 163),
  (x => 168, y => 163),
  (x => 169, y => 163),
  (x => 170, y => 163),
  (x => 187, y => 163),
  (x => 188, y => 163),
  (x => 189, y => 163),
  (x => 190, y => 163),
  (x => 191, y => 163),
  (x => 192, y => 163),
  (x => 193, y => 163),
  (x => 201, y => 163),
  (x => 202, y => 163),
  (x => 203, y => 163),
  (x => 204, y => 163),
  (x => 205, y => 163),
  (x => 206, y => 163),
  (x => 217, y => 163),
  (x => 218, y => 163),
  (x => 219, y => 163),
  (x => 220, y => 163),
  (x => 221, y => 163),
  (x => 222, y => 163),
  (x => 231, y => 163),
  (x => 232, y => 163),
  (x => 233, y => 163),
  (x => 234, y => 163),
  (x => 235, y => 163),
  (x => 236, y => 163),
  (x => 237, y => 163),
  (x => 248, y => 163),
  (x => 249, y => 163),
  (x => 250, y => 163),
  (x => 251, y => 163),
  (x => 252, y => 163),
  (x => 253, y => 163),
  (x => 254, y => 163),
  (x => 266, y => 163),
  (x => 267, y => 163),
  (x => 268, y => 163),
  (x => 269, y => 163),
  (x => 270, y => 163),
  (x => 271, y => 163),
  (x => 272, y => 163),
  (x => 279, y => 163),
  (x => 280, y => 163),
  (x => 281, y => 163),
  (x => 282, y => 163),
  (x => 283, y => 163),
  (x => 284, y => 163),
  (x => 285, y => 163),
  (x => 324, y => 163),
  (x => 325, y => 163),
  (x => 326, y => 163),
  (x => 327, y => 163),
  (x => 328, y => 163),
  (x => 329, y => 163),
  (x => 330, y => 163),
  (x => 331, y => 163),
  (x => 350, y => 163),
  (x => 351, y => 163),
  (x => 352, y => 163),
  (x => 353, y => 163),
  (x => 354, y => 163),
  (x => 355, y => 163),
  (x => 356, y => 163),
  (x => 357, y => 163),
  (x => 368, y => 163),
  (x => 369, y => 163),
  (x => 370, y => 163),
  (x => 371, y => 163),
  (x => 372, y => 163),
  (x => 373, y => 163),
  (x => 378, y => 163),
  (x => 379, y => 163),
  (x => 380, y => 163),
  (x => 381, y => 163),
  (x => 382, y => 163),
  (x => 383, y => 163),
  (x => 394, y => 163),
  (x => 395, y => 163),
  (x => 396, y => 163),
  (x => 397, y => 163),
  (x => 398, y => 163),
  (x => 399, y => 163),
  (x => 424, y => 163),
  (x => 425, y => 163),
  (x => 426, y => 163),
  (x => 427, y => 163),
  (x => 428, y => 163),
  (x => 429, y => 163),
  (x => 430, y => 163),
  (x => 163, y => 164),
  (x => 164, y => 164),
  (x => 165, y => 164),
  (x => 166, y => 164),
  (x => 167, y => 164),
  (x => 168, y => 164),
  (x => 169, y => 164),
  (x => 170, y => 164),
  (x => 171, y => 164),
  (x => 187, y => 164),
  (x => 188, y => 164),
  (x => 189, y => 164),
  (x => 190, y => 164),
  (x => 191, y => 164),
  (x => 192, y => 164),
  (x => 193, y => 164),
  (x => 200, y => 164),
  (x => 201, y => 164),
  (x => 202, y => 164),
  (x => 203, y => 164),
  (x => 204, y => 164),
  (x => 205, y => 164),
  (x => 206, y => 164),
  (x => 217, y => 164),
  (x => 218, y => 164),
  (x => 219, y => 164),
  (x => 220, y => 164),
  (x => 221, y => 164),
  (x => 222, y => 164),
  (x => 231, y => 164),
  (x => 232, y => 164),
  (x => 233, y => 164),
  (x => 234, y => 164),
  (x => 235, y => 164),
  (x => 236, y => 164),
  (x => 237, y => 164),
  (x => 248, y => 164),
  (x => 249, y => 164),
  (x => 250, y => 164),
  (x => 251, y => 164),
  (x => 252, y => 164),
  (x => 253, y => 164),
  (x => 254, y => 164),
  (x => 266, y => 164),
  (x => 267, y => 164),
  (x => 268, y => 164),
  (x => 269, y => 164),
  (x => 270, y => 164),
  (x => 271, y => 164),
  (x => 272, y => 164),
  (x => 279, y => 164),
  (x => 280, y => 164),
  (x => 281, y => 164),
  (x => 282, y => 164),
  (x => 283, y => 164),
  (x => 284, y => 164),
  (x => 285, y => 164),
  (x => 325, y => 164),
  (x => 326, y => 164),
  (x => 327, y => 164),
  (x => 328, y => 164),
  (x => 329, y => 164),
  (x => 330, y => 164),
  (x => 331, y => 164),
  (x => 332, y => 164),
  (x => 349, y => 164),
  (x => 350, y => 164),
  (x => 351, y => 164),
  (x => 352, y => 164),
  (x => 353, y => 164),
  (x => 354, y => 164),
  (x => 355, y => 164),
  (x => 356, y => 164),
  (x => 368, y => 164),
  (x => 369, y => 164),
  (x => 370, y => 164),
  (x => 371, y => 164),
  (x => 372, y => 164),
  (x => 373, y => 164),
  (x => 378, y => 164),
  (x => 379, y => 164),
  (x => 380, y => 164),
  (x => 381, y => 164),
  (x => 382, y => 164),
  (x => 383, y => 164),
  (x => 394, y => 164),
  (x => 395, y => 164),
  (x => 396, y => 164),
  (x => 397, y => 164),
  (x => 398, y => 164),
  (x => 399, y => 164),
  (x => 424, y => 164),
  (x => 425, y => 164),
  (x => 426, y => 164),
  (x => 427, y => 164),
  (x => 428, y => 164),
  (x => 429, y => 164),
  (x => 430, y => 164),
  (x => 164, y => 165),
  (x => 165, y => 165),
  (x => 166, y => 165),
  (x => 167, y => 165),
  (x => 168, y => 165),
  (x => 169, y => 165),
  (x => 170, y => 165),
  (x => 171, y => 165),
  (x => 172, y => 165),
  (x => 187, y => 165),
  (x => 188, y => 165),
  (x => 189, y => 165),
  (x => 190, y => 165),
  (x => 191, y => 165),
  (x => 192, y => 165),
  (x => 193, y => 165),
  (x => 200, y => 165),
  (x => 201, y => 165),
  (x => 202, y => 165),
  (x => 203, y => 165),
  (x => 204, y => 165),
  (x => 205, y => 165),
  (x => 217, y => 165),
  (x => 218, y => 165),
  (x => 219, y => 165),
  (x => 220, y => 165),
  (x => 221, y => 165),
  (x => 222, y => 165),
  (x => 231, y => 165),
  (x => 232, y => 165),
  (x => 233, y => 165),
  (x => 234, y => 165),
  (x => 235, y => 165),
  (x => 236, y => 165),
  (x => 237, y => 165),
  (x => 248, y => 165),
  (x => 249, y => 165),
  (x => 250, y => 165),
  (x => 251, y => 165),
  (x => 252, y => 165),
  (x => 253, y => 165),
  (x => 254, y => 165),
  (x => 266, y => 165),
  (x => 267, y => 165),
  (x => 268, y => 165),
  (x => 269, y => 165),
  (x => 270, y => 165),
  (x => 271, y => 165),
  (x => 272, y => 165),
  (x => 279, y => 165),
  (x => 280, y => 165),
  (x => 281, y => 165),
  (x => 282, y => 165),
  (x => 283, y => 165),
  (x => 284, y => 165),
  (x => 285, y => 165),
  (x => 325, y => 165),
  (x => 326, y => 165),
  (x => 327, y => 165),
  (x => 328, y => 165),
  (x => 329, y => 165),
  (x => 330, y => 165),
  (x => 331, y => 165),
  (x => 332, y => 165),
  (x => 349, y => 165),
  (x => 350, y => 165),
  (x => 351, y => 165),
  (x => 352, y => 165),
  (x => 353, y => 165),
  (x => 354, y => 165),
  (x => 355, y => 165),
  (x => 356, y => 165),
  (x => 369, y => 165),
  (x => 370, y => 165),
  (x => 371, y => 165),
  (x => 372, y => 165),
  (x => 373, y => 165),
  (x => 374, y => 165),
  (x => 378, y => 165),
  (x => 379, y => 165),
  (x => 380, y => 165),
  (x => 381, y => 165),
  (x => 382, y => 165),
  (x => 383, y => 165),
  (x => 394, y => 165),
  (x => 395, y => 165),
  (x => 396, y => 165),
  (x => 397, y => 165),
  (x => 398, y => 165),
  (x => 399, y => 165),
  (x => 424, y => 165),
  (x => 425, y => 165),
  (x => 426, y => 165),
  (x => 427, y => 165),
  (x => 428, y => 165),
  (x => 429, y => 165),
  (x => 430, y => 165),
  (x => 164, y => 166),
  (x => 165, y => 166),
  (x => 166, y => 166),
  (x => 167, y => 166),
  (x => 168, y => 166),
  (x => 169, y => 166),
  (x => 170, y => 166),
  (x => 171, y => 166),
  (x => 172, y => 166),
  (x => 187, y => 166),
  (x => 188, y => 166),
  (x => 189, y => 166),
  (x => 190, y => 166),
  (x => 191, y => 166),
  (x => 192, y => 166),
  (x => 193, y => 166),
  (x => 200, y => 166),
  (x => 201, y => 166),
  (x => 202, y => 166),
  (x => 203, y => 166),
  (x => 204, y => 166),
  (x => 205, y => 166),
  (x => 216, y => 166),
  (x => 217, y => 166),
  (x => 218, y => 166),
  (x => 219, y => 166),
  (x => 220, y => 166),
  (x => 221, y => 166),
  (x => 222, y => 166),
  (x => 231, y => 166),
  (x => 232, y => 166),
  (x => 233, y => 166),
  (x => 234, y => 166),
  (x => 235, y => 166),
  (x => 236, y => 166),
  (x => 237, y => 166),
  (x => 248, y => 166),
  (x => 249, y => 166),
  (x => 250, y => 166),
  (x => 251, y => 166),
  (x => 252, y => 166),
  (x => 253, y => 166),
  (x => 254, y => 166),
  (x => 266, y => 166),
  (x => 267, y => 166),
  (x => 268, y => 166),
  (x => 269, y => 166),
  (x => 270, y => 166),
  (x => 271, y => 166),
  (x => 272, y => 166),
  (x => 279, y => 166),
  (x => 280, y => 166),
  (x => 281, y => 166),
  (x => 282, y => 166),
  (x => 283, y => 166),
  (x => 284, y => 166),
  (x => 285, y => 166),
  (x => 325, y => 166),
  (x => 326, y => 166),
  (x => 327, y => 166),
  (x => 328, y => 166),
  (x => 329, y => 166),
  (x => 330, y => 166),
  (x => 331, y => 166),
  (x => 332, y => 166),
  (x => 333, y => 166),
  (x => 348, y => 166),
  (x => 349, y => 166),
  (x => 350, y => 166),
  (x => 351, y => 166),
  (x => 352, y => 166),
  (x => 353, y => 166),
  (x => 354, y => 166),
  (x => 355, y => 166),
  (x => 356, y => 166),
  (x => 369, y => 166),
  (x => 370, y => 166),
  (x => 371, y => 166),
  (x => 372, y => 166),
  (x => 373, y => 166),
  (x => 374, y => 166),
  (x => 378, y => 166),
  (x => 379, y => 166),
  (x => 380, y => 166),
  (x => 381, y => 166),
  (x => 382, y => 166),
  (x => 394, y => 166),
  (x => 395, y => 166),
  (x => 396, y => 166),
  (x => 397, y => 166),
  (x => 398, y => 166),
  (x => 399, y => 166),
  (x => 400, y => 166),
  (x => 424, y => 166),
  (x => 425, y => 166),
  (x => 426, y => 166),
  (x => 427, y => 166),
  (x => 428, y => 166),
  (x => 429, y => 166),
  (x => 430, y => 166),
  (x => 165, y => 167),
  (x => 166, y => 167),
  (x => 167, y => 167),
  (x => 168, y => 167),
  (x => 169, y => 167),
  (x => 170, y => 167),
  (x => 171, y => 167),
  (x => 172, y => 167),
  (x => 173, y => 167),
  (x => 187, y => 167),
  (x => 188, y => 167),
  (x => 189, y => 167),
  (x => 190, y => 167),
  (x => 191, y => 167),
  (x => 192, y => 167),
  (x => 193, y => 167),
  (x => 200, y => 167),
  (x => 201, y => 167),
  (x => 202, y => 167),
  (x => 203, y => 167),
  (x => 204, y => 167),
  (x => 205, y => 167),
  (x => 216, y => 167),
  (x => 217, y => 167),
  (x => 218, y => 167),
  (x => 219, y => 167),
  (x => 220, y => 167),
  (x => 221, y => 167),
  (x => 222, y => 167),
  (x => 231, y => 167),
  (x => 232, y => 167),
  (x => 233, y => 167),
  (x => 234, y => 167),
  (x => 235, y => 167),
  (x => 236, y => 167),
  (x => 237, y => 167),
  (x => 248, y => 167),
  (x => 249, y => 167),
  (x => 250, y => 167),
  (x => 251, y => 167),
  (x => 252, y => 167),
  (x => 253, y => 167),
  (x => 254, y => 167),
  (x => 266, y => 167),
  (x => 267, y => 167),
  (x => 268, y => 167),
  (x => 269, y => 167),
  (x => 270, y => 167),
  (x => 271, y => 167),
  (x => 272, y => 167),
  (x => 280, y => 167),
  (x => 281, y => 167),
  (x => 282, y => 167),
  (x => 283, y => 167),
  (x => 284, y => 167),
  (x => 285, y => 167),
  (x => 326, y => 167),
  (x => 327, y => 167),
  (x => 328, y => 167),
  (x => 329, y => 167),
  (x => 330, y => 167),
  (x => 331, y => 167),
  (x => 332, y => 167),
  (x => 333, y => 167),
  (x => 334, y => 167),
  (x => 347, y => 167),
  (x => 348, y => 167),
  (x => 349, y => 167),
  (x => 350, y => 167),
  (x => 351, y => 167),
  (x => 352, y => 167),
  (x => 353, y => 167),
  (x => 354, y => 167),
  (x => 355, y => 167),
  (x => 369, y => 167),
  (x => 370, y => 167),
  (x => 371, y => 167),
  (x => 372, y => 167),
  (x => 373, y => 167),
  (x => 374, y => 167),
  (x => 377, y => 167),
  (x => 378, y => 167),
  (x => 379, y => 167),
  (x => 380, y => 167),
  (x => 381, y => 167),
  (x => 382, y => 167),
  (x => 394, y => 167),
  (x => 395, y => 167),
  (x => 396, y => 167),
  (x => 397, y => 167),
  (x => 398, y => 167),
  (x => 399, y => 167),
  (x => 400, y => 167),
  (x => 424, y => 167),
  (x => 425, y => 167),
  (x => 426, y => 167),
  (x => 427, y => 167),
  (x => 428, y => 167),
  (x => 429, y => 167),
  (x => 430, y => 167),
  (x => 165, y => 168),
  (x => 166, y => 168),
  (x => 167, y => 168),
  (x => 168, y => 168),
  (x => 169, y => 168),
  (x => 170, y => 168),
  (x => 171, y => 168),
  (x => 172, y => 168),
  (x => 173, y => 168),
  (x => 174, y => 168),
  (x => 187, y => 168),
  (x => 188, y => 168),
  (x => 189, y => 168),
  (x => 190, y => 168),
  (x => 191, y => 168),
  (x => 192, y => 168),
  (x => 193, y => 168),
  (x => 200, y => 168),
  (x => 201, y => 168),
  (x => 202, y => 168),
  (x => 203, y => 168),
  (x => 204, y => 168),
  (x => 205, y => 168),
  (x => 216, y => 168),
  (x => 217, y => 168),
  (x => 218, y => 168),
  (x => 219, y => 168),
  (x => 220, y => 168),
  (x => 221, y => 168),
  (x => 222, y => 168),
  (x => 231, y => 168),
  (x => 232, y => 168),
  (x => 233, y => 168),
  (x => 234, y => 168),
  (x => 235, y => 168),
  (x => 236, y => 168),
  (x => 237, y => 168),
  (x => 248, y => 168),
  (x => 249, y => 168),
  (x => 250, y => 168),
  (x => 251, y => 168),
  (x => 252, y => 168),
  (x => 253, y => 168),
  (x => 254, y => 168),
  (x => 266, y => 168),
  (x => 267, y => 168),
  (x => 268, y => 168),
  (x => 269, y => 168),
  (x => 270, y => 168),
  (x => 271, y => 168),
  (x => 272, y => 168),
  (x => 280, y => 168),
  (x => 281, y => 168),
  (x => 282, y => 168),
  (x => 283, y => 168),
  (x => 284, y => 168),
  (x => 285, y => 168),
  (x => 286, y => 168),
  (x => 326, y => 168),
  (x => 327, y => 168),
  (x => 328, y => 168),
  (x => 329, y => 168),
  (x => 330, y => 168),
  (x => 331, y => 168),
  (x => 332, y => 168),
  (x => 333, y => 168),
  (x => 334, y => 168),
  (x => 335, y => 168),
  (x => 346, y => 168),
  (x => 347, y => 168),
  (x => 348, y => 168),
  (x => 349, y => 168),
  (x => 350, y => 168),
  (x => 351, y => 168),
  (x => 352, y => 168),
  (x => 353, y => 168),
  (x => 354, y => 168),
  (x => 355, y => 168),
  (x => 369, y => 168),
  (x => 370, y => 168),
  (x => 371, y => 168),
  (x => 372, y => 168),
  (x => 373, y => 168),
  (x => 374, y => 168),
  (x => 377, y => 168),
  (x => 378, y => 168),
  (x => 379, y => 168),
  (x => 380, y => 168),
  (x => 381, y => 168),
  (x => 382, y => 168),
  (x => 394, y => 168),
  (x => 395, y => 168),
  (x => 396, y => 168),
  (x => 397, y => 168),
  (x => 398, y => 168),
  (x => 399, y => 168),
  (x => 400, y => 168),
  (x => 424, y => 168),
  (x => 425, y => 168),
  (x => 426, y => 168),
  (x => 427, y => 168),
  (x => 428, y => 168),
  (x => 429, y => 168),
  (x => 430, y => 168),
  (x => 165, y => 169),
  (x => 166, y => 169),
  (x => 167, y => 169),
  (x => 168, y => 169),
  (x => 169, y => 169),
  (x => 170, y => 169),
  (x => 171, y => 169),
  (x => 172, y => 169),
  (x => 173, y => 169),
  (x => 174, y => 169),
  (x => 175, y => 169),
  (x => 176, y => 169),
  (x => 187, y => 169),
  (x => 188, y => 169),
  (x => 189, y => 169),
  (x => 190, y => 169),
  (x => 191, y => 169),
  (x => 192, y => 169),
  (x => 193, y => 169),
  (x => 200, y => 169),
  (x => 201, y => 169),
  (x => 202, y => 169),
  (x => 203, y => 169),
  (x => 204, y => 169),
  (x => 205, y => 169),
  (x => 206, y => 169),
  (x => 215, y => 169),
  (x => 216, y => 169),
  (x => 217, y => 169),
  (x => 218, y => 169),
  (x => 219, y => 169),
  (x => 220, y => 169),
  (x => 221, y => 169),
  (x => 222, y => 169),
  (x => 231, y => 169),
  (x => 232, y => 169),
  (x => 233, y => 169),
  (x => 234, y => 169),
  (x => 235, y => 169),
  (x => 236, y => 169),
  (x => 237, y => 169),
  (x => 248, y => 169),
  (x => 249, y => 169),
  (x => 250, y => 169),
  (x => 251, y => 169),
  (x => 252, y => 169),
  (x => 253, y => 169),
  (x => 254, y => 169),
  (x => 266, y => 169),
  (x => 267, y => 169),
  (x => 268, y => 169),
  (x => 269, y => 169),
  (x => 270, y => 169),
  (x => 271, y => 169),
  (x => 272, y => 169),
  (x => 280, y => 169),
  (x => 281, y => 169),
  (x => 282, y => 169),
  (x => 283, y => 169),
  (x => 284, y => 169),
  (x => 285, y => 169),
  (x => 286, y => 169),
  (x => 327, y => 169),
  (x => 328, y => 169),
  (x => 329, y => 169),
  (x => 330, y => 169),
  (x => 331, y => 169),
  (x => 332, y => 169),
  (x => 333, y => 169),
  (x => 334, y => 169),
  (x => 335, y => 169),
  (x => 336, y => 169),
  (x => 345, y => 169),
  (x => 346, y => 169),
  (x => 347, y => 169),
  (x => 348, y => 169),
  (x => 349, y => 169),
  (x => 350, y => 169),
  (x => 351, y => 169),
  (x => 352, y => 169),
  (x => 353, y => 169),
  (x => 354, y => 169),
  (x => 370, y => 169),
  (x => 371, y => 169),
  (x => 372, y => 169),
  (x => 373, y => 169),
  (x => 374, y => 169),
  (x => 377, y => 169),
  (x => 378, y => 169),
  (x => 379, y => 169),
  (x => 380, y => 169),
  (x => 381, y => 169),
  (x => 395, y => 169),
  (x => 396, y => 169),
  (x => 397, y => 169),
  (x => 398, y => 169),
  (x => 399, y => 169),
  (x => 400, y => 169),
  (x => 401, y => 169),
  (x => 424, y => 169),
  (x => 425, y => 169),
  (x => 426, y => 169),
  (x => 427, y => 169),
  (x => 428, y => 169),
  (x => 429, y => 169),
  (x => 430, y => 169),
  (x => 166, y => 170),
  (x => 167, y => 170),
  (x => 168, y => 170),
  (x => 169, y => 170),
  (x => 170, y => 170),
  (x => 171, y => 170),
  (x => 172, y => 170),
  (x => 173, y => 170),
  (x => 174, y => 170),
  (x => 175, y => 170),
  (x => 176, y => 170),
  (x => 177, y => 170),
  (x => 178, y => 170),
  (x => 184, y => 170),
  (x => 185, y => 170),
  (x => 186, y => 170),
  (x => 187, y => 170),
  (x => 188, y => 170),
  (x => 189, y => 170),
  (x => 190, y => 170),
  (x => 191, y => 170),
  (x => 192, y => 170),
  (x => 193, y => 170),
  (x => 200, y => 170),
  (x => 201, y => 170),
  (x => 202, y => 170),
  (x => 203, y => 170),
  (x => 204, y => 170),
  (x => 205, y => 170),
  (x => 206, y => 170),
  (x => 214, y => 170),
  (x => 215, y => 170),
  (x => 216, y => 170),
  (x => 217, y => 170),
  (x => 218, y => 170),
  (x => 219, y => 170),
  (x => 220, y => 170),
  (x => 221, y => 170),
  (x => 222, y => 170),
  (x => 231, y => 170),
  (x => 232, y => 170),
  (x => 233, y => 170),
  (x => 234, y => 170),
  (x => 235, y => 170),
  (x => 236, y => 170),
  (x => 237, y => 170),
  (x => 248, y => 170),
  (x => 249, y => 170),
  (x => 250, y => 170),
  (x => 251, y => 170),
  (x => 252, y => 170),
  (x => 253, y => 170),
  (x => 254, y => 170),
  (x => 266, y => 170),
  (x => 267, y => 170),
  (x => 268, y => 170),
  (x => 269, y => 170),
  (x => 270, y => 170),
  (x => 271, y => 170),
  (x => 272, y => 170),
  (x => 280, y => 170),
  (x => 281, y => 170),
  (x => 282, y => 170),
  (x => 283, y => 170),
  (x => 284, y => 170),
  (x => 285, y => 170),
  (x => 286, y => 170),
  (x => 287, y => 170),
  (x => 327, y => 170),
  (x => 328, y => 170),
  (x => 329, y => 170),
  (x => 330, y => 170),
  (x => 331, y => 170),
  (x => 332, y => 170),
  (x => 333, y => 170),
  (x => 334, y => 170),
  (x => 335, y => 170),
  (x => 336, y => 170),
  (x => 337, y => 170),
  (x => 338, y => 170),
  (x => 339, y => 170),
  (x => 340, y => 170),
  (x => 341, y => 170),
  (x => 342, y => 170),
  (x => 343, y => 170),
  (x => 344, y => 170),
  (x => 345, y => 170),
  (x => 346, y => 170),
  (x => 347, y => 170),
  (x => 348, y => 170),
  (x => 349, y => 170),
  (x => 350, y => 170),
  (x => 351, y => 170),
  (x => 352, y => 170),
  (x => 353, y => 170),
  (x => 354, y => 170),
  (x => 370, y => 170),
  (x => 371, y => 170),
  (x => 372, y => 170),
  (x => 373, y => 170),
  (x => 374, y => 170),
  (x => 377, y => 170),
  (x => 378, y => 170),
  (x => 379, y => 170),
  (x => 380, y => 170),
  (x => 381, y => 170),
  (x => 395, y => 170),
  (x => 396, y => 170),
  (x => 397, y => 170),
  (x => 398, y => 170),
  (x => 399, y => 170),
  (x => 400, y => 170),
  (x => 401, y => 170),
  (x => 402, y => 170),
  (x => 415, y => 170),
  (x => 424, y => 170),
  (x => 425, y => 170),
  (x => 426, y => 170),
  (x => 427, y => 170),
  (x => 428, y => 170),
  (x => 429, y => 170),
  (x => 430, y => 170),
  (x => 167, y => 171),
  (x => 168, y => 171),
  (x => 169, y => 171),
  (x => 170, y => 171),
  (x => 171, y => 171),
  (x => 172, y => 171),
  (x => 173, y => 171),
  (x => 174, y => 171),
  (x => 175, y => 171),
  (x => 176, y => 171),
  (x => 177, y => 171),
  (x => 178, y => 171),
  (x => 179, y => 171),
  (x => 180, y => 171),
  (x => 181, y => 171),
  (x => 182, y => 171),
  (x => 183, y => 171),
  (x => 184, y => 171),
  (x => 185, y => 171),
  (x => 186, y => 171),
  (x => 187, y => 171),
  (x => 188, y => 171),
  (x => 189, y => 171),
  (x => 190, y => 171),
  (x => 191, y => 171),
  (x => 192, y => 171),
  (x => 193, y => 171),
  (x => 200, y => 171),
  (x => 201, y => 171),
  (x => 202, y => 171),
  (x => 203, y => 171),
  (x => 204, y => 171),
  (x => 205, y => 171),
  (x => 206, y => 171),
  (x => 207, y => 171),
  (x => 213, y => 171),
  (x => 214, y => 171),
  (x => 215, y => 171),
  (x => 216, y => 171),
  (x => 217, y => 171),
  (x => 218, y => 171),
  (x => 219, y => 171),
  (x => 220, y => 171),
  (x => 221, y => 171),
  (x => 222, y => 171),
  (x => 231, y => 171),
  (x => 232, y => 171),
  (x => 233, y => 171),
  (x => 234, y => 171),
  (x => 235, y => 171),
  (x => 236, y => 171),
  (x => 237, y => 171),
  (x => 248, y => 171),
  (x => 249, y => 171),
  (x => 250, y => 171),
  (x => 251, y => 171),
  (x => 252, y => 171),
  (x => 253, y => 171),
  (x => 254, y => 171),
  (x => 266, y => 171),
  (x => 267, y => 171),
  (x => 268, y => 171),
  (x => 269, y => 171),
  (x => 270, y => 171),
  (x => 271, y => 171),
  (x => 272, y => 171),
  (x => 281, y => 171),
  (x => 282, y => 171),
  (x => 283, y => 171),
  (x => 284, y => 171),
  (x => 285, y => 171),
  (x => 286, y => 171),
  (x => 287, y => 171),
  (x => 288, y => 171),
  (x => 289, y => 171),
  (x => 299, y => 171),
  (x => 300, y => 171),
  (x => 328, y => 171),
  (x => 329, y => 171),
  (x => 330, y => 171),
  (x => 331, y => 171),
  (x => 332, y => 171),
  (x => 333, y => 171),
  (x => 334, y => 171),
  (x => 335, y => 171),
  (x => 336, y => 171),
  (x => 337, y => 171),
  (x => 338, y => 171),
  (x => 339, y => 171),
  (x => 340, y => 171),
  (x => 341, y => 171),
  (x => 342, y => 171),
  (x => 343, y => 171),
  (x => 344, y => 171),
  (x => 345, y => 171),
  (x => 346, y => 171),
  (x => 347, y => 171),
  (x => 348, y => 171),
  (x => 349, y => 171),
  (x => 350, y => 171),
  (x => 351, y => 171),
  (x => 352, y => 171),
  (x => 353, y => 171),
  (x => 370, y => 171),
  (x => 371, y => 171),
  (x => 372, y => 171),
  (x => 373, y => 171),
  (x => 374, y => 171),
  (x => 375, y => 171),
  (x => 376, y => 171),
  (x => 377, y => 171),
  (x => 378, y => 171),
  (x => 379, y => 171),
  (x => 380, y => 171),
  (x => 381, y => 171),
  (x => 395, y => 171),
  (x => 396, y => 171),
  (x => 397, y => 171),
  (x => 398, y => 171),
  (x => 399, y => 171),
  (x => 400, y => 171),
  (x => 401, y => 171),
  (x => 402, y => 171),
  (x => 403, y => 171),
  (x => 413, y => 171),
  (x => 414, y => 171),
  (x => 415, y => 171),
  (x => 424, y => 171),
  (x => 425, y => 171),
  (x => 426, y => 171),
  (x => 427, y => 171),
  (x => 428, y => 171),
  (x => 429, y => 171),
  (x => 430, y => 171),
  (x => 167, y => 172),
  (x => 168, y => 172),
  (x => 169, y => 172),
  (x => 170, y => 172),
  (x => 171, y => 172),
  (x => 172, y => 172),
  (x => 173, y => 172),
  (x => 174, y => 172),
  (x => 175, y => 172),
  (x => 176, y => 172),
  (x => 177, y => 172),
  (x => 178, y => 172),
  (x => 179, y => 172),
  (x => 180, y => 172),
  (x => 181, y => 172),
  (x => 182, y => 172),
  (x => 183, y => 172),
  (x => 184, y => 172),
  (x => 185, y => 172),
  (x => 186, y => 172),
  (x => 187, y => 172),
  (x => 188, y => 172),
  (x => 189, y => 172),
  (x => 190, y => 172),
  (x => 191, y => 172),
  (x => 192, y => 172),
  (x => 193, y => 172),
  (x => 200, y => 172),
  (x => 201, y => 172),
  (x => 202, y => 172),
  (x => 203, y => 172),
  (x => 204, y => 172),
  (x => 205, y => 172),
  (x => 206, y => 172),
  (x => 207, y => 172),
  (x => 208, y => 172),
  (x => 209, y => 172),
  (x => 210, y => 172),
  (x => 211, y => 172),
  (x => 212, y => 172),
  (x => 213, y => 172),
  (x => 214, y => 172),
  (x => 215, y => 172),
  (x => 216, y => 172),
  (x => 217, y => 172),
  (x => 218, y => 172),
  (x => 219, y => 172),
  (x => 220, y => 172),
  (x => 221, y => 172),
  (x => 222, y => 172),
  (x => 231, y => 172),
  (x => 232, y => 172),
  (x => 233, y => 172),
  (x => 234, y => 172),
  (x => 235, y => 172),
  (x => 236, y => 172),
  (x => 237, y => 172),
  (x => 248, y => 172),
  (x => 249, y => 172),
  (x => 250, y => 172),
  (x => 251, y => 172),
  (x => 252, y => 172),
  (x => 253, y => 172),
  (x => 254, y => 172),
  (x => 266, y => 172),
  (x => 267, y => 172),
  (x => 268, y => 172),
  (x => 269, y => 172),
  (x => 270, y => 172),
  (x => 271, y => 172),
  (x => 272, y => 172),
  (x => 281, y => 172),
  (x => 282, y => 172),
  (x => 283, y => 172),
  (x => 284, y => 172),
  (x => 285, y => 172),
  (x => 286, y => 172),
  (x => 287, y => 172),
  (x => 288, y => 172),
  (x => 289, y => 172),
  (x => 290, y => 172),
  (x => 291, y => 172),
  (x => 292, y => 172),
  (x => 293, y => 172),
  (x => 294, y => 172),
  (x => 295, y => 172),
  (x => 296, y => 172),
  (x => 297, y => 172),
  (x => 298, y => 172),
  (x => 299, y => 172),
  (x => 300, y => 172),
  (x => 329, y => 172),
  (x => 330, y => 172),
  (x => 331, y => 172),
  (x => 332, y => 172),
  (x => 333, y => 172),
  (x => 334, y => 172),
  (x => 335, y => 172),
  (x => 336, y => 172),
  (x => 337, y => 172),
  (x => 338, y => 172),
  (x => 339, y => 172),
  (x => 340, y => 172),
  (x => 341, y => 172),
  (x => 342, y => 172),
  (x => 343, y => 172),
  (x => 344, y => 172),
  (x => 345, y => 172),
  (x => 346, y => 172),
  (x => 347, y => 172),
  (x => 348, y => 172),
  (x => 349, y => 172),
  (x => 350, y => 172),
  (x => 351, y => 172),
  (x => 352, y => 172),
  (x => 370, y => 172),
  (x => 371, y => 172),
  (x => 372, y => 172),
  (x => 373, y => 172),
  (x => 374, y => 172),
  (x => 375, y => 172),
  (x => 376, y => 172),
  (x => 377, y => 172),
  (x => 378, y => 172),
  (x => 379, y => 172),
  (x => 380, y => 172),
  (x => 381, y => 172),
  (x => 396, y => 172),
  (x => 397, y => 172),
  (x => 398, y => 172),
  (x => 399, y => 172),
  (x => 400, y => 172),
  (x => 401, y => 172),
  (x => 402, y => 172),
  (x => 403, y => 172),
  (x => 404, y => 172),
  (x => 405, y => 172),
  (x => 406, y => 172),
  (x => 407, y => 172),
  (x => 408, y => 172),
  (x => 409, y => 172),
  (x => 410, y => 172),
  (x => 411, y => 172),
  (x => 412, y => 172),
  (x => 413, y => 172),
  (x => 414, y => 172),
  (x => 415, y => 172),
  (x => 424, y => 172),
  (x => 425, y => 172),
  (x => 426, y => 172),
  (x => 427, y => 172),
  (x => 428, y => 172),
  (x => 429, y => 172),
  (x => 430, y => 172),
  (x => 168, y => 173),
  (x => 169, y => 173),
  (x => 170, y => 173),
  (x => 171, y => 173),
  (x => 172, y => 173),
  (x => 173, y => 173),
  (x => 174, y => 173),
  (x => 175, y => 173),
  (x => 176, y => 173),
  (x => 177, y => 173),
  (x => 178, y => 173),
  (x => 179, y => 173),
  (x => 180, y => 173),
  (x => 181, y => 173),
  (x => 182, y => 173),
  (x => 183, y => 173),
  (x => 184, y => 173),
  (x => 185, y => 173),
  (x => 186, y => 173),
  (x => 187, y => 173),
  (x => 188, y => 173),
  (x => 189, y => 173),
  (x => 190, y => 173),
  (x => 191, y => 173),
  (x => 192, y => 173),
  (x => 193, y => 173),
  (x => 201, y => 173),
  (x => 202, y => 173),
  (x => 203, y => 173),
  (x => 204, y => 173),
  (x => 205, y => 173),
  (x => 206, y => 173),
  (x => 207, y => 173),
  (x => 208, y => 173),
  (x => 209, y => 173),
  (x => 210, y => 173),
  (x => 211, y => 173),
  (x => 212, y => 173),
  (x => 213, y => 173),
  (x => 214, y => 173),
  (x => 217, y => 173),
  (x => 218, y => 173),
  (x => 219, y => 173),
  (x => 220, y => 173),
  (x => 221, y => 173),
  (x => 222, y => 173),
  (x => 231, y => 173),
  (x => 232, y => 173),
  (x => 233, y => 173),
  (x => 234, y => 173),
  (x => 235, y => 173),
  (x => 236, y => 173),
  (x => 237, y => 173),
  (x => 248, y => 173),
  (x => 249, y => 173),
  (x => 250, y => 173),
  (x => 251, y => 173),
  (x => 252, y => 173),
  (x => 253, y => 173),
  (x => 254, y => 173),
  (x => 266, y => 173),
  (x => 267, y => 173),
  (x => 268, y => 173),
  (x => 269, y => 173),
  (x => 270, y => 173),
  (x => 271, y => 173),
  (x => 272, y => 173),
  (x => 282, y => 173),
  (x => 283, y => 173),
  (x => 284, y => 173),
  (x => 285, y => 173),
  (x => 286, y => 173),
  (x => 287, y => 173),
  (x => 288, y => 173),
  (x => 289, y => 173),
  (x => 290, y => 173),
  (x => 291, y => 173),
  (x => 292, y => 173),
  (x => 293, y => 173),
  (x => 294, y => 173),
  (x => 295, y => 173),
  (x => 296, y => 173),
  (x => 297, y => 173),
  (x => 298, y => 173),
  (x => 299, y => 173),
  (x => 300, y => 173),
  (x => 329, y => 173),
  (x => 330, y => 173),
  (x => 331, y => 173),
  (x => 332, y => 173),
  (x => 333, y => 173),
  (x => 334, y => 173),
  (x => 335, y => 173),
  (x => 336, y => 173),
  (x => 337, y => 173),
  (x => 338, y => 173),
  (x => 339, y => 173),
  (x => 340, y => 173),
  (x => 341, y => 173),
  (x => 342, y => 173),
  (x => 343, y => 173),
  (x => 344, y => 173),
  (x => 345, y => 173),
  (x => 346, y => 173),
  (x => 347, y => 173),
  (x => 348, y => 173),
  (x => 349, y => 173),
  (x => 350, y => 173),
  (x => 351, y => 173),
  (x => 371, y => 173),
  (x => 372, y => 173),
  (x => 373, y => 173),
  (x => 374, y => 173),
  (x => 375, y => 173),
  (x => 376, y => 173),
  (x => 377, y => 173),
  (x => 378, y => 173),
  (x => 379, y => 173),
  (x => 380, y => 173),
  (x => 396, y => 173),
  (x => 397, y => 173),
  (x => 398, y => 173),
  (x => 399, y => 173),
  (x => 400, y => 173),
  (x => 401, y => 173),
  (x => 402, y => 173),
  (x => 403, y => 173),
  (x => 404, y => 173),
  (x => 405, y => 173),
  (x => 406, y => 173),
  (x => 407, y => 173),
  (x => 408, y => 173),
  (x => 409, y => 173),
  (x => 410, y => 173),
  (x => 411, y => 173),
  (x => 412, y => 173),
  (x => 413, y => 173),
  (x => 414, y => 173),
  (x => 415, y => 173),
  (x => 424, y => 173),
  (x => 425, y => 173),
  (x => 426, y => 173),
  (x => 427, y => 173),
  (x => 428, y => 173),
  (x => 429, y => 173),
  (x => 430, y => 173),
  (x => 169, y => 174),
  (x => 170, y => 174),
  (x => 171, y => 174),
  (x => 172, y => 174),
  (x => 173, y => 174),
  (x => 174, y => 174),
  (x => 175, y => 174),
  (x => 176, y => 174),
  (x => 177, y => 174),
  (x => 178, y => 174),
  (x => 179, y => 174),
  (x => 180, y => 174),
  (x => 181, y => 174),
  (x => 182, y => 174),
  (x => 183, y => 174),
  (x => 184, y => 174),
  (x => 185, y => 174),
  (x => 186, y => 174),
  (x => 187, y => 174),
  (x => 188, y => 174),
  (x => 189, y => 174),
  (x => 190, y => 174),
  (x => 191, y => 174),
  (x => 192, y => 174),
  (x => 193, y => 174),
  (x => 201, y => 174),
  (x => 202, y => 174),
  (x => 203, y => 174),
  (x => 204, y => 174),
  (x => 205, y => 174),
  (x => 206, y => 174),
  (x => 207, y => 174),
  (x => 208, y => 174),
  (x => 209, y => 174),
  (x => 210, y => 174),
  (x => 211, y => 174),
  (x => 212, y => 174),
  (x => 213, y => 174),
  (x => 217, y => 174),
  (x => 218, y => 174),
  (x => 219, y => 174),
  (x => 220, y => 174),
  (x => 221, y => 174),
  (x => 222, y => 174),
  (x => 231, y => 174),
  (x => 232, y => 174),
  (x => 233, y => 174),
  (x => 234, y => 174),
  (x => 235, y => 174),
  (x => 236, y => 174),
  (x => 237, y => 174),
  (x => 248, y => 174),
  (x => 249, y => 174),
  (x => 250, y => 174),
  (x => 251, y => 174),
  (x => 252, y => 174),
  (x => 253, y => 174),
  (x => 254, y => 174),
  (x => 266, y => 174),
  (x => 267, y => 174),
  (x => 268, y => 174),
  (x => 269, y => 174),
  (x => 270, y => 174),
  (x => 271, y => 174),
  (x => 272, y => 174),
  (x => 283, y => 174),
  (x => 284, y => 174),
  (x => 285, y => 174),
  (x => 286, y => 174),
  (x => 287, y => 174),
  (x => 288, y => 174),
  (x => 289, y => 174),
  (x => 290, y => 174),
  (x => 291, y => 174),
  (x => 292, y => 174),
  (x => 293, y => 174),
  (x => 294, y => 174),
  (x => 295, y => 174),
  (x => 296, y => 174),
  (x => 297, y => 174),
  (x => 298, y => 174),
  (x => 299, y => 174),
  (x => 300, y => 174),
  (x => 330, y => 174),
  (x => 331, y => 174),
  (x => 332, y => 174),
  (x => 333, y => 174),
  (x => 334, y => 174),
  (x => 335, y => 174),
  (x => 336, y => 174),
  (x => 337, y => 174),
  (x => 338, y => 174),
  (x => 339, y => 174),
  (x => 340, y => 174),
  (x => 341, y => 174),
  (x => 342, y => 174),
  (x => 343, y => 174),
  (x => 344, y => 174),
  (x => 345, y => 174),
  (x => 346, y => 174),
  (x => 347, y => 174),
  (x => 348, y => 174),
  (x => 349, y => 174),
  (x => 350, y => 174),
  (x => 351, y => 174),
  (x => 371, y => 174),
  (x => 372, y => 174),
  (x => 373, y => 174),
  (x => 374, y => 174),
  (x => 375, y => 174),
  (x => 376, y => 174),
  (x => 377, y => 174),
  (x => 378, y => 174),
  (x => 379, y => 174),
  (x => 380, y => 174),
  (x => 397, y => 174),
  (x => 398, y => 174),
  (x => 399, y => 174),
  (x => 400, y => 174),
  (x => 401, y => 174),
  (x => 402, y => 174),
  (x => 403, y => 174),
  (x => 404, y => 174),
  (x => 405, y => 174),
  (x => 406, y => 174),
  (x => 407, y => 174),
  (x => 408, y => 174),
  (x => 409, y => 174),
  (x => 410, y => 174),
  (x => 411, y => 174),
  (x => 412, y => 174),
  (x => 413, y => 174),
  (x => 414, y => 174),
  (x => 415, y => 174),
  (x => 424, y => 174),
  (x => 425, y => 174),
  (x => 426, y => 174),
  (x => 427, y => 174),
  (x => 428, y => 174),
  (x => 429, y => 174),
  (x => 430, y => 174),
  (x => 171, y => 175),
  (x => 172, y => 175),
  (x => 173, y => 175),
  (x => 174, y => 175),
  (x => 175, y => 175),
  (x => 176, y => 175),
  (x => 177, y => 175),
  (x => 178, y => 175),
  (x => 179, y => 175),
  (x => 180, y => 175),
  (x => 181, y => 175),
  (x => 182, y => 175),
  (x => 183, y => 175),
  (x => 184, y => 175),
  (x => 185, y => 175),
  (x => 186, y => 175),
  (x => 187, y => 175),
  (x => 188, y => 175),
  (x => 189, y => 175),
  (x => 190, y => 175),
  (x => 191, y => 175),
  (x => 192, y => 175),
  (x => 202, y => 175),
  (x => 203, y => 175),
  (x => 204, y => 175),
  (x => 205, y => 175),
  (x => 206, y => 175),
  (x => 207, y => 175),
  (x => 208, y => 175),
  (x => 209, y => 175),
  (x => 210, y => 175),
  (x => 211, y => 175),
  (x => 212, y => 175),
  (x => 213, y => 175),
  (x => 217, y => 175),
  (x => 218, y => 175),
  (x => 219, y => 175),
  (x => 220, y => 175),
  (x => 221, y => 175),
  (x => 222, y => 175),
  (x => 231, y => 175),
  (x => 232, y => 175),
  (x => 233, y => 175),
  (x => 234, y => 175),
  (x => 235, y => 175),
  (x => 236, y => 175),
  (x => 237, y => 175),
  (x => 248, y => 175),
  (x => 249, y => 175),
  (x => 250, y => 175),
  (x => 251, y => 175),
  (x => 252, y => 175),
  (x => 253, y => 175),
  (x => 254, y => 175),
  (x => 266, y => 175),
  (x => 267, y => 175),
  (x => 268, y => 175),
  (x => 269, y => 175),
  (x => 270, y => 175),
  (x => 271, y => 175),
  (x => 272, y => 175),
  (x => 283, y => 175),
  (x => 284, y => 175),
  (x => 285, y => 175),
  (x => 286, y => 175),
  (x => 287, y => 175),
  (x => 288, y => 175),
  (x => 289, y => 175),
  (x => 290, y => 175),
  (x => 291, y => 175),
  (x => 292, y => 175),
  (x => 293, y => 175),
  (x => 294, y => 175),
  (x => 295, y => 175),
  (x => 296, y => 175),
  (x => 297, y => 175),
  (x => 298, y => 175),
  (x => 299, y => 175),
  (x => 300, y => 175),
  (x => 331, y => 175),
  (x => 332, y => 175),
  (x => 333, y => 175),
  (x => 334, y => 175),
  (x => 335, y => 175),
  (x => 336, y => 175),
  (x => 337, y => 175),
  (x => 338, y => 175),
  (x => 339, y => 175),
  (x => 340, y => 175),
  (x => 341, y => 175),
  (x => 342, y => 175),
  (x => 343, y => 175),
  (x => 344, y => 175),
  (x => 345, y => 175),
  (x => 346, y => 175),
  (x => 347, y => 175),
  (x => 348, y => 175),
  (x => 349, y => 175),
  (x => 371, y => 175),
  (x => 372, y => 175),
  (x => 373, y => 175),
  (x => 374, y => 175),
  (x => 375, y => 175),
  (x => 376, y => 175),
  (x => 377, y => 175),
  (x => 378, y => 175),
  (x => 379, y => 175),
  (x => 380, y => 175),
  (x => 398, y => 175),
  (x => 399, y => 175),
  (x => 400, y => 175),
  (x => 401, y => 175),
  (x => 402, y => 175),
  (x => 403, y => 175),
  (x => 404, y => 175),
  (x => 405, y => 175),
  (x => 406, y => 175),
  (x => 407, y => 175),
  (x => 408, y => 175),
  (x => 409, y => 175),
  (x => 410, y => 175),
  (x => 411, y => 175),
  (x => 412, y => 175),
  (x => 413, y => 175),
  (x => 414, y => 175),
  (x => 415, y => 175),
  (x => 424, y => 175),
  (x => 425, y => 175),
  (x => 426, y => 175),
  (x => 427, y => 175),
  (x => 428, y => 175),
  (x => 429, y => 175),
  (x => 430, y => 175),
  (x => 172, y => 176),
  (x => 173, y => 176),
  (x => 174, y => 176),
  (x => 175, y => 176),
  (x => 176, y => 176),
  (x => 177, y => 176),
  (x => 178, y => 176),
  (x => 179, y => 176),
  (x => 180, y => 176),
  (x => 181, y => 176),
  (x => 182, y => 176),
  (x => 183, y => 176),
  (x => 184, y => 176),
  (x => 185, y => 176),
  (x => 186, y => 176),
  (x => 187, y => 176),
  (x => 188, y => 176),
  (x => 189, y => 176),
  (x => 190, y => 176),
  (x => 202, y => 176),
  (x => 203, y => 176),
  (x => 204, y => 176),
  (x => 205, y => 176),
  (x => 206, y => 176),
  (x => 207, y => 176),
  (x => 208, y => 176),
  (x => 209, y => 176),
  (x => 210, y => 176),
  (x => 211, y => 176),
  (x => 212, y => 176),
  (x => 217, y => 176),
  (x => 218, y => 176),
  (x => 219, y => 176),
  (x => 220, y => 176),
  (x => 221, y => 176),
  (x => 222, y => 176),
  (x => 231, y => 176),
  (x => 232, y => 176),
  (x => 233, y => 176),
  (x => 234, y => 176),
  (x => 235, y => 176),
  (x => 236, y => 176),
  (x => 237, y => 176),
  (x => 248, y => 176),
  (x => 249, y => 176),
  (x => 250, y => 176),
  (x => 251, y => 176),
  (x => 252, y => 176),
  (x => 253, y => 176),
  (x => 254, y => 176),
  (x => 266, y => 176),
  (x => 267, y => 176),
  (x => 268, y => 176),
  (x => 269, y => 176),
  (x => 270, y => 176),
  (x => 271, y => 176),
  (x => 272, y => 176),
  (x => 285, y => 176),
  (x => 286, y => 176),
  (x => 287, y => 176),
  (x => 288, y => 176),
  (x => 289, y => 176),
  (x => 290, y => 176),
  (x => 291, y => 176),
  (x => 292, y => 176),
  (x => 293, y => 176),
  (x => 294, y => 176),
  (x => 295, y => 176),
  (x => 296, y => 176),
  (x => 297, y => 176),
  (x => 298, y => 176),
  (x => 299, y => 176),
  (x => 300, y => 176),
  (x => 333, y => 176),
  (x => 334, y => 176),
  (x => 335, y => 176),
  (x => 336, y => 176),
  (x => 337, y => 176),
  (x => 338, y => 176),
  (x => 339, y => 176),
  (x => 340, y => 176),
  (x => 341, y => 176),
  (x => 342, y => 176),
  (x => 343, y => 176),
  (x => 344, y => 176),
  (x => 345, y => 176),
  (x => 346, y => 176),
  (x => 347, y => 176),
  (x => 348, y => 176),
  (x => 371, y => 176),
  (x => 372, y => 176),
  (x => 373, y => 176),
  (x => 374, y => 176),
  (x => 375, y => 176),
  (x => 376, y => 176),
  (x => 377, y => 176),
  (x => 378, y => 176),
  (x => 379, y => 176),
  (x => 399, y => 176),
  (x => 400, y => 176),
  (x => 401, y => 176),
  (x => 402, y => 176),
  (x => 403, y => 176),
  (x => 404, y => 176),
  (x => 405, y => 176),
  (x => 406, y => 176),
  (x => 407, y => 176),
  (x => 408, y => 176),
  (x => 409, y => 176),
  (x => 410, y => 176),
  (x => 411, y => 176),
  (x => 412, y => 176),
  (x => 413, y => 176),
  (x => 414, y => 176),
  (x => 424, y => 176),
  (x => 425, y => 176),
  (x => 426, y => 176),
  (x => 427, y => 176),
  (x => 428, y => 176),
  (x => 429, y => 176),
  (x => 430, y => 176),
  (x => 174, y => 177),
  (x => 175, y => 177),
  (x => 176, y => 177),
  (x => 177, y => 177),
  (x => 178, y => 177),
  (x => 179, y => 177),
  (x => 180, y => 177),
  (x => 181, y => 177),
  (x => 182, y => 177),
  (x => 183, y => 177),
  (x => 184, y => 177),
  (x => 185, y => 177),
  (x => 186, y => 177),
  (x => 187, y => 177),
  (x => 188, y => 177),
  (x => 204, y => 177),
  (x => 205, y => 177),
  (x => 206, y => 177),
  (x => 207, y => 177),
  (x => 208, y => 177),
  (x => 209, y => 177),
  (x => 210, y => 177),
  (x => 211, y => 177),
  (x => 216, y => 177),
  (x => 217, y => 177),
  (x => 218, y => 177),
  (x => 219, y => 177),
  (x => 220, y => 177),
  (x => 221, y => 177),
  (x => 222, y => 177),
  (x => 231, y => 177),
  (x => 232, y => 177),
  (x => 233, y => 177),
  (x => 234, y => 177),
  (x => 235, y => 177),
  (x => 236, y => 177),
  (x => 237, y => 177),
  (x => 248, y => 177),
  (x => 249, y => 177),
  (x => 250, y => 177),
  (x => 251, y => 177),
  (x => 252, y => 177),
  (x => 253, y => 177),
  (x => 254, y => 177),
  (x => 265, y => 177),
  (x => 266, y => 177),
  (x => 267, y => 177),
  (x => 268, y => 177),
  (x => 269, y => 177),
  (x => 270, y => 177),
  (x => 271, y => 177),
  (x => 272, y => 177),
  (x => 286, y => 177),
  (x => 287, y => 177),
  (x => 288, y => 177),
  (x => 289, y => 177),
  (x => 290, y => 177),
  (x => 291, y => 177),
  (x => 292, y => 177),
  (x => 293, y => 177),
  (x => 294, y => 177),
  (x => 295, y => 177),
  (x => 296, y => 177),
  (x => 297, y => 177),
  (x => 298, y => 177),
  (x => 335, y => 177),
  (x => 336, y => 177),
  (x => 337, y => 177),
  (x => 338, y => 177),
  (x => 339, y => 177),
  (x => 340, y => 177),
  (x => 341, y => 177),
  (x => 342, y => 177),
  (x => 343, y => 177),
  (x => 344, y => 177),
  (x => 345, y => 177),
  (x => 346, y => 177),
  (x => 372, y => 177),
  (x => 373, y => 177),
  (x => 374, y => 177),
  (x => 375, y => 177),
  (x => 376, y => 177),
  (x => 377, y => 177),
  (x => 378, y => 177),
  (x => 379, y => 177),
  (x => 401, y => 177),
  (x => 402, y => 177),
  (x => 403, y => 177),
  (x => 404, y => 177),
  (x => 405, y => 177),
  (x => 406, y => 177),
  (x => 407, y => 177),
  (x => 408, y => 177),
  (x => 409, y => 177),
  (x => 410, y => 177),
  (x => 411, y => 177),
  (x => 412, y => 177),
  (x => 424, y => 177),
  (x => 425, y => 177),
  (x => 426, y => 177),
  (x => 427, y => 177),
  (x => 428, y => 177),
  (x => 429, y => 177),
  (x => 430, y => 177),
  (x => 178, y => 178),
  (x => 179, y => 178),
  (x => 180, y => 178),
  (x => 181, y => 178),
  (x => 182, y => 178),
  (x => 183, y => 178),
  (x => 206, y => 178),
  (x => 207, y => 178),
  (x => 208, y => 178),
  (x => 290, y => 178),
  (x => 291, y => 178),
  (x => 292, y => 178),
  (x => 293, y => 178),
  (x => 294, y => 178),
  (x => 338, y => 178),
  (x => 339, y => 178),
  (x => 340, y => 178),
  (x => 341, y => 178),
  (x => 342, y => 178),
  (x => 404, y => 178),
  (x => 405, y => 178),
  (x => 406, y => 178),
  (x => 407, y => 178),
  (x => 408, y => 178),
  (x => 409, y => 178),
  (x => 228, y => 222),
  (x => 229, y => 222),
  (x => 230, y => 222),
  (x => 231, y => 222),
  (x => 368, y => 222),
  (x => 369, y => 222),
  (x => 209, y => 223),
  (x => 210, y => 223),
  (x => 211, y => 223),
  (x => 212, y => 223),
  (x => 213, y => 223),
  (x => 214, y => 223),
  (x => 215, y => 223),
  (x => 216, y => 223),
  (x => 217, y => 223),
  (x => 228, y => 223),
  (x => 229, y => 223),
  (x => 230, y => 223),
  (x => 231, y => 223),
  (x => 334, y => 223),
  (x => 335, y => 223),
  (x => 336, y => 223),
  (x => 337, y => 223),
  (x => 347, y => 223),
  (x => 348, y => 223),
  (x => 349, y => 223),
  (x => 350, y => 223),
  (x => 360, y => 223),
  (x => 361, y => 223),
  (x => 362, y => 223),
  (x => 367, y => 223),
  (x => 368, y => 223),
  (x => 369, y => 223),
  (x => 370, y => 223),
  (x => 209, y => 224),
  (x => 210, y => 224),
  (x => 211, y => 224),
  (x => 212, y => 224),
  (x => 213, y => 224),
  (x => 214, y => 224),
  (x => 215, y => 224),
  (x => 216, y => 224),
  (x => 217, y => 224),
  (x => 218, y => 224),
  (x => 219, y => 224),
  (x => 220, y => 224),
  (x => 228, y => 224),
  (x => 229, y => 224),
  (x => 230, y => 224),
  (x => 231, y => 224),
  (x => 313, y => 224),
  (x => 314, y => 224),
  (x => 315, y => 224),
  (x => 316, y => 224),
  (x => 317, y => 224),
  (x => 318, y => 224),
  (x => 334, y => 224),
  (x => 335, y => 224),
  (x => 336, y => 224),
  (x => 337, y => 224),
  (x => 347, y => 224),
  (x => 348, y => 224),
  (x => 349, y => 224),
  (x => 350, y => 224),
  (x => 360, y => 224),
  (x => 361, y => 224),
  (x => 362, y => 224),
  (x => 367, y => 224),
  (x => 368, y => 224),
  (x => 369, y => 224),
  (x => 370, y => 224),
  (x => 209, y => 225),
  (x => 210, y => 225),
  (x => 211, y => 225),
  (x => 212, y => 225),
  (x => 213, y => 225),
  (x => 214, y => 225),
  (x => 215, y => 225),
  (x => 216, y => 225),
  (x => 217, y => 225),
  (x => 218, y => 225),
  (x => 219, y => 225),
  (x => 220, y => 225),
  (x => 221, y => 225),
  (x => 228, y => 225),
  (x => 229, y => 225),
  (x => 230, y => 225),
  (x => 231, y => 225),
  (x => 312, y => 225),
  (x => 313, y => 225),
  (x => 314, y => 225),
  (x => 315, y => 225),
  (x => 316, y => 225),
  (x => 317, y => 225),
  (x => 318, y => 225),
  (x => 319, y => 225),
  (x => 320, y => 225),
  (x => 335, y => 225),
  (x => 336, y => 225),
  (x => 337, y => 225),
  (x => 347, y => 225),
  (x => 348, y => 225),
  (x => 349, y => 225),
  (x => 350, y => 225),
  (x => 351, y => 225),
  (x => 360, y => 225),
  (x => 361, y => 225),
  (x => 362, y => 225),
  (x => 367, y => 225),
  (x => 368, y => 225),
  (x => 369, y => 225),
  (x => 370, y => 225),
  (x => 209, y => 226),
  (x => 210, y => 226),
  (x => 211, y => 226),
  (x => 212, y => 226),
  (x => 213, y => 226),
  (x => 214, y => 226),
  (x => 215, y => 226),
  (x => 216, y => 226),
  (x => 217, y => 226),
  (x => 218, y => 226),
  (x => 219, y => 226),
  (x => 220, y => 226),
  (x => 221, y => 226),
  (x => 222, y => 226),
  (x => 228, y => 226),
  (x => 229, y => 226),
  (x => 230, y => 226),
  (x => 231, y => 226),
  (x => 311, y => 226),
  (x => 312, y => 226),
  (x => 313, y => 226),
  (x => 314, y => 226),
  (x => 315, y => 226),
  (x => 316, y => 226),
  (x => 317, y => 226),
  (x => 318, y => 226),
  (x => 319, y => 226),
  (x => 320, y => 226),
  (x => 321, y => 226),
  (x => 335, y => 226),
  (x => 336, y => 226),
  (x => 337, y => 226),
  (x => 347, y => 226),
  (x => 348, y => 226),
  (x => 349, y => 226),
  (x => 350, y => 226),
  (x => 351, y => 226),
  (x => 359, y => 226),
  (x => 360, y => 226),
  (x => 361, y => 226),
  (x => 362, y => 226),
  (x => 368, y => 226),
  (x => 369, y => 226),
  (x => 209, y => 227),
  (x => 210, y => 227),
  (x => 211, y => 227),
  (x => 212, y => 227),
  (x => 217, y => 227),
  (x => 218, y => 227),
  (x => 219, y => 227),
  (x => 220, y => 227),
  (x => 221, y => 227),
  (x => 222, y => 227),
  (x => 228, y => 227),
  (x => 229, y => 227),
  (x => 230, y => 227),
  (x => 231, y => 227),
  (x => 311, y => 227),
  (x => 312, y => 227),
  (x => 313, y => 227),
  (x => 314, y => 227),
  (x => 315, y => 227),
  (x => 316, y => 227),
  (x => 317, y => 227),
  (x => 318, y => 227),
  (x => 319, y => 227),
  (x => 320, y => 227),
  (x => 321, y => 227),
  (x => 335, y => 227),
  (x => 336, y => 227),
  (x => 337, y => 227),
  (x => 338, y => 227),
  (x => 346, y => 227),
  (x => 347, y => 227),
  (x => 348, y => 227),
  (x => 349, y => 227),
  (x => 350, y => 227),
  (x => 351, y => 227),
  (x => 359, y => 227),
  (x => 360, y => 227),
  (x => 361, y => 227),
  (x => 362, y => 227),
  (x => 209, y => 228),
  (x => 210, y => 228),
  (x => 211, y => 228),
  (x => 212, y => 228),
  (x => 219, y => 228),
  (x => 220, y => 228),
  (x => 221, y => 228),
  (x => 222, y => 228),
  (x => 223, y => 228),
  (x => 228, y => 228),
  (x => 229, y => 228),
  (x => 230, y => 228),
  (x => 231, y => 228),
  (x => 311, y => 228),
  (x => 312, y => 228),
  (x => 318, y => 228),
  (x => 319, y => 228),
  (x => 320, y => 228),
  (x => 321, y => 228),
  (x => 322, y => 228),
  (x => 335, y => 228),
  (x => 336, y => 228),
  (x => 337, y => 228),
  (x => 338, y => 228),
  (x => 346, y => 228),
  (x => 347, y => 228),
  (x => 348, y => 228),
  (x => 349, y => 228),
  (x => 350, y => 228),
  (x => 351, y => 228),
  (x => 359, y => 228),
  (x => 360, y => 228),
  (x => 361, y => 228),
  (x => 209, y => 229),
  (x => 210, y => 229),
  (x => 211, y => 229),
  (x => 212, y => 229),
  (x => 220, y => 229),
  (x => 221, y => 229),
  (x => 222, y => 229),
  (x => 223, y => 229),
  (x => 228, y => 229),
  (x => 229, y => 229),
  (x => 230, y => 229),
  (x => 231, y => 229),
  (x => 319, y => 229),
  (x => 320, y => 229),
  (x => 321, y => 229),
  (x => 322, y => 229),
  (x => 335, y => 229),
  (x => 336, y => 229),
  (x => 337, y => 229),
  (x => 338, y => 229),
  (x => 346, y => 229),
  (x => 347, y => 229),
  (x => 348, y => 229),
  (x => 349, y => 229),
  (x => 350, y => 229),
  (x => 351, y => 229),
  (x => 359, y => 229),
  (x => 360, y => 229),
  (x => 361, y => 229),
  (x => 209, y => 230),
  (x => 210, y => 230),
  (x => 211, y => 230),
  (x => 212, y => 230),
  (x => 220, y => 230),
  (x => 221, y => 230),
  (x => 222, y => 230),
  (x => 223, y => 230),
  (x => 228, y => 230),
  (x => 229, y => 230),
  (x => 230, y => 230),
  (x => 231, y => 230),
  (x => 319, y => 230),
  (x => 320, y => 230),
  (x => 321, y => 230),
  (x => 322, y => 230),
  (x => 335, y => 230),
  (x => 336, y => 230),
  (x => 337, y => 230),
  (x => 338, y => 230),
  (x => 346, y => 230),
  (x => 347, y => 230),
  (x => 350, y => 230),
  (x => 351, y => 230),
  (x => 352, y => 230),
  (x => 359, y => 230),
  (x => 360, y => 230),
  (x => 361, y => 230),
  (x => 209, y => 231),
  (x => 210, y => 231),
  (x => 211, y => 231),
  (x => 212, y => 231),
  (x => 220, y => 231),
  (x => 221, y => 231),
  (x => 222, y => 231),
  (x => 223, y => 231),
  (x => 228, y => 231),
  (x => 229, y => 231),
  (x => 230, y => 231),
  (x => 231, y => 231),
  (x => 242, y => 231),
  (x => 243, y => 231),
  (x => 276, y => 231),
  (x => 277, y => 231),
  (x => 296, y => 231),
  (x => 319, y => 231),
  (x => 320, y => 231),
  (x => 321, y => 231),
  (x => 322, y => 231),
  (x => 336, y => 231),
  (x => 337, y => 231),
  (x => 338, y => 231),
  (x => 346, y => 231),
  (x => 347, y => 231),
  (x => 350, y => 231),
  (x => 351, y => 231),
  (x => 352, y => 231),
  (x => 359, y => 231),
  (x => 360, y => 231),
  (x => 361, y => 231),
  (x => 385, y => 231),
  (x => 386, y => 231),
  (x => 399, y => 231),
  (x => 400, y => 231),
  (x => 401, y => 231),
  (x => 209, y => 232),
  (x => 210, y => 232),
  (x => 211, y => 232),
  (x => 212, y => 232),
  (x => 220, y => 232),
  (x => 221, y => 232),
  (x => 222, y => 232),
  (x => 223, y => 232),
  (x => 228, y => 232),
  (x => 229, y => 232),
  (x => 230, y => 232),
  (x => 231, y => 232),
  (x => 238, y => 232),
  (x => 239, y => 232),
  (x => 240, y => 232),
  (x => 241, y => 232),
  (x => 242, y => 232),
  (x => 243, y => 232),
  (x => 244, y => 232),
  (x => 245, y => 232),
  (x => 246, y => 232),
  (x => 252, y => 232),
  (x => 253, y => 232),
  (x => 254, y => 232),
  (x => 255, y => 232),
  (x => 264, y => 232),
  (x => 265, y => 232),
  (x => 266, y => 232),
  (x => 267, y => 232),
  (x => 274, y => 232),
  (x => 275, y => 232),
  (x => 276, y => 232),
  (x => 277, y => 232),
  (x => 278, y => 232),
  (x => 279, y => 232),
  (x => 280, y => 232),
  (x => 288, y => 232),
  (x => 289, y => 232),
  (x => 290, y => 232),
  (x => 291, y => 232),
  (x => 294, y => 232),
  (x => 295, y => 232),
  (x => 296, y => 232),
  (x => 319, y => 232),
  (x => 320, y => 232),
  (x => 321, y => 232),
  (x => 322, y => 232),
  (x => 336, y => 232),
  (x => 337, y => 232),
  (x => 338, y => 232),
  (x => 345, y => 232),
  (x => 346, y => 232),
  (x => 347, y => 232),
  (x => 350, y => 232),
  (x => 351, y => 232),
  (x => 352, y => 232),
  (x => 358, y => 232),
  (x => 359, y => 232),
  (x => 360, y => 232),
  (x => 361, y => 232),
  (x => 367, y => 232),
  (x => 368, y => 232),
  (x => 369, y => 232),
  (x => 370, y => 232),
  (x => 376, y => 232),
  (x => 377, y => 232),
  (x => 378, y => 232),
  (x => 379, y => 232),
  (x => 383, y => 232),
  (x => 384, y => 232),
  (x => 385, y => 232),
  (x => 386, y => 232),
  (x => 387, y => 232),
  (x => 397, y => 232),
  (x => 398, y => 232),
  (x => 399, y => 232),
  (x => 400, y => 232),
  (x => 401, y => 232),
  (x => 402, y => 232),
  (x => 403, y => 232),
  (x => 209, y => 233),
  (x => 210, y => 233),
  (x => 211, y => 233),
  (x => 212, y => 233),
  (x => 220, y => 233),
  (x => 221, y => 233),
  (x => 222, y => 233),
  (x => 223, y => 233),
  (x => 228, y => 233),
  (x => 229, y => 233),
  (x => 230, y => 233),
  (x => 231, y => 233),
  (x => 238, y => 233),
  (x => 239, y => 233),
  (x => 240, y => 233),
  (x => 241, y => 233),
  (x => 242, y => 233),
  (x => 243, y => 233),
  (x => 244, y => 233),
  (x => 245, y => 233),
  (x => 246, y => 233),
  (x => 247, y => 233),
  (x => 253, y => 233),
  (x => 254, y => 233),
  (x => 255, y => 233),
  (x => 256, y => 233),
  (x => 264, y => 233),
  (x => 265, y => 233),
  (x => 266, y => 233),
  (x => 273, y => 233),
  (x => 274, y => 233),
  (x => 275, y => 233),
  (x => 276, y => 233),
  (x => 277, y => 233),
  (x => 278, y => 233),
  (x => 279, y => 233),
  (x => 280, y => 233),
  (x => 281, y => 233),
  (x => 288, y => 233),
  (x => 289, y => 233),
  (x => 290, y => 233),
  (x => 294, y => 233),
  (x => 295, y => 233),
  (x => 296, y => 233),
  (x => 319, y => 233),
  (x => 320, y => 233),
  (x => 321, y => 233),
  (x => 322, y => 233),
  (x => 336, y => 233),
  (x => 337, y => 233),
  (x => 338, y => 233),
  (x => 339, y => 233),
  (x => 345, y => 233),
  (x => 346, y => 233),
  (x => 347, y => 233),
  (x => 350, y => 233),
  (x => 351, y => 233),
  (x => 352, y => 233),
  (x => 358, y => 233),
  (x => 359, y => 233),
  (x => 360, y => 233),
  (x => 367, y => 233),
  (x => 368, y => 233),
  (x => 369, y => 233),
  (x => 370, y => 233),
  (x => 376, y => 233),
  (x => 377, y => 233),
  (x => 378, y => 233),
  (x => 379, y => 233),
  (x => 382, y => 233),
  (x => 383, y => 233),
  (x => 384, y => 233),
  (x => 385, y => 233),
  (x => 386, y => 233),
  (x => 387, y => 233),
  (x => 388, y => 233),
  (x => 396, y => 233),
  (x => 397, y => 233),
  (x => 398, y => 233),
  (x => 399, y => 233),
  (x => 400, y => 233),
  (x => 401, y => 233),
  (x => 402, y => 233),
  (x => 403, y => 233),
  (x => 209, y => 234),
  (x => 210, y => 234),
  (x => 211, y => 234),
  (x => 212, y => 234),
  (x => 220, y => 234),
  (x => 221, y => 234),
  (x => 222, y => 234),
  (x => 223, y => 234),
  (x => 228, y => 234),
  (x => 229, y => 234),
  (x => 230, y => 234),
  (x => 231, y => 234),
  (x => 238, y => 234),
  (x => 239, y => 234),
  (x => 240, y => 234),
  (x => 241, y => 234),
  (x => 243, y => 234),
  (x => 244, y => 234),
  (x => 245, y => 234),
  (x => 246, y => 234),
  (x => 247, y => 234),
  (x => 253, y => 234),
  (x => 254, y => 234),
  (x => 255, y => 234),
  (x => 256, y => 234),
  (x => 264, y => 234),
  (x => 265, y => 234),
  (x => 266, y => 234),
  (x => 272, y => 234),
  (x => 273, y => 234),
  (x => 274, y => 234),
  (x => 275, y => 234),
  (x => 276, y => 234),
  (x => 278, y => 234),
  (x => 279, y => 234),
  (x => 280, y => 234),
  (x => 281, y => 234),
  (x => 288, y => 234),
  (x => 289, y => 234),
  (x => 290, y => 234),
  (x => 293, y => 234),
  (x => 294, y => 234),
  (x => 295, y => 234),
  (x => 296, y => 234),
  (x => 319, y => 234),
  (x => 320, y => 234),
  (x => 321, y => 234),
  (x => 322, y => 234),
  (x => 336, y => 234),
  (x => 337, y => 234),
  (x => 338, y => 234),
  (x => 339, y => 234),
  (x => 345, y => 234),
  (x => 346, y => 234),
  (x => 350, y => 234),
  (x => 351, y => 234),
  (x => 352, y => 234),
  (x => 358, y => 234),
  (x => 359, y => 234),
  (x => 360, y => 234),
  (x => 367, y => 234),
  (x => 368, y => 234),
  (x => 369, y => 234),
  (x => 370, y => 234),
  (x => 376, y => 234),
  (x => 377, y => 234),
  (x => 378, y => 234),
  (x => 379, y => 234),
  (x => 382, y => 234),
  (x => 383, y => 234),
  (x => 384, y => 234),
  (x => 385, y => 234),
  (x => 386, y => 234),
  (x => 387, y => 234),
  (x => 388, y => 234),
  (x => 389, y => 234),
  (x => 395, y => 234),
  (x => 396, y => 234),
  (x => 397, y => 234),
  (x => 398, y => 234),
  (x => 399, y => 234),
  (x => 400, y => 234),
  (x => 401, y => 234),
  (x => 402, y => 234),
  (x => 403, y => 234),
  (x => 209, y => 235),
  (x => 210, y => 235),
  (x => 211, y => 235),
  (x => 212, y => 235),
  (x => 220, y => 235),
  (x => 221, y => 235),
  (x => 222, y => 235),
  (x => 223, y => 235),
  (x => 228, y => 235),
  (x => 229, y => 235),
  (x => 230, y => 235),
  (x => 231, y => 235),
  (x => 238, y => 235),
  (x => 245, y => 235),
  (x => 246, y => 235),
  (x => 247, y => 235),
  (x => 254, y => 235),
  (x => 255, y => 235),
  (x => 256, y => 235),
  (x => 264, y => 235),
  (x => 265, y => 235),
  (x => 266, y => 235),
  (x => 272, y => 235),
  (x => 273, y => 235),
  (x => 274, y => 235),
  (x => 280, y => 235),
  (x => 281, y => 235),
  (x => 282, y => 235),
  (x => 288, y => 235),
  (x => 289, y => 235),
  (x => 290, y => 235),
  (x => 291, y => 235),
  (x => 292, y => 235),
  (x => 293, y => 235),
  (x => 294, y => 235),
  (x => 295, y => 235),
  (x => 296, y => 235),
  (x => 319, y => 235),
  (x => 320, y => 235),
  (x => 321, y => 235),
  (x => 337, y => 235),
  (x => 338, y => 235),
  (x => 339, y => 235),
  (x => 345, y => 235),
  (x => 346, y => 235),
  (x => 350, y => 235),
  (x => 351, y => 235),
  (x => 352, y => 235),
  (x => 358, y => 235),
  (x => 359, y => 235),
  (x => 360, y => 235),
  (x => 367, y => 235),
  (x => 368, y => 235),
  (x => 369, y => 235),
  (x => 370, y => 235),
  (x => 376, y => 235),
  (x => 377, y => 235),
  (x => 378, y => 235),
  (x => 379, y => 235),
  (x => 380, y => 235),
  (x => 381, y => 235),
  (x => 385, y => 235),
  (x => 386, y => 235),
  (x => 387, y => 235),
  (x => 388, y => 235),
  (x => 389, y => 235),
  (x => 395, y => 235),
  (x => 396, y => 235),
  (x => 397, y => 235),
  (x => 209, y => 236),
  (x => 210, y => 236),
  (x => 211, y => 236),
  (x => 212, y => 236),
  (x => 219, y => 236),
  (x => 220, y => 236),
  (x => 221, y => 236),
  (x => 222, y => 236),
  (x => 228, y => 236),
  (x => 229, y => 236),
  (x => 230, y => 236),
  (x => 231, y => 236),
  (x => 246, y => 236),
  (x => 247, y => 236),
  (x => 248, y => 236),
  (x => 254, y => 236),
  (x => 255, y => 236),
  (x => 256, y => 236),
  (x => 263, y => 236),
  (x => 264, y => 236),
  (x => 265, y => 236),
  (x => 271, y => 236),
  (x => 272, y => 236),
  (x => 273, y => 236),
  (x => 280, y => 236),
  (x => 281, y => 236),
  (x => 282, y => 236),
  (x => 288, y => 236),
  (x => 289, y => 236),
  (x => 290, y => 236),
  (x => 291, y => 236),
  (x => 292, y => 236),
  (x => 318, y => 236),
  (x => 319, y => 236),
  (x => 320, y => 236),
  (x => 321, y => 236),
  (x => 337, y => 236),
  (x => 338, y => 236),
  (x => 339, y => 236),
  (x => 345, y => 236),
  (x => 346, y => 236),
  (x => 351, y => 236),
  (x => 352, y => 236),
  (x => 353, y => 236),
  (x => 358, y => 236),
  (x => 359, y => 236),
  (x => 360, y => 236),
  (x => 367, y => 236),
  (x => 368, y => 236),
  (x => 369, y => 236),
  (x => 370, y => 236),
  (x => 376, y => 236),
  (x => 377, y => 236),
  (x => 378, y => 236),
  (x => 379, y => 236),
  (x => 380, y => 236),
  (x => 386, y => 236),
  (x => 387, y => 236),
  (x => 388, y => 236),
  (x => 389, y => 236),
  (x => 394, y => 236),
  (x => 395, y => 236),
  (x => 396, y => 236),
  (x => 397, y => 236),
  (x => 209, y => 237),
  (x => 210, y => 237),
  (x => 211, y => 237),
  (x => 212, y => 237),
  (x => 218, y => 237),
  (x => 219, y => 237),
  (x => 220, y => 237),
  (x => 221, y => 237),
  (x => 222, y => 237),
  (x => 228, y => 237),
  (x => 229, y => 237),
  (x => 230, y => 237),
  (x => 231, y => 237),
  (x => 246, y => 237),
  (x => 247, y => 237),
  (x => 248, y => 237),
  (x => 254, y => 237),
  (x => 255, y => 237),
  (x => 256, y => 237),
  (x => 263, y => 237),
  (x => 264, y => 237),
  (x => 265, y => 237),
  (x => 271, y => 237),
  (x => 272, y => 237),
  (x => 273, y => 237),
  (x => 281, y => 237),
  (x => 282, y => 237),
  (x => 288, y => 237),
  (x => 289, y => 237),
  (x => 290, y => 237),
  (x => 291, y => 237),
  (x => 318, y => 237),
  (x => 319, y => 237),
  (x => 320, y => 237),
  (x => 321, y => 237),
  (x => 337, y => 237),
  (x => 338, y => 237),
  (x => 339, y => 237),
  (x => 344, y => 237),
  (x => 345, y => 237),
  (x => 346, y => 237),
  (x => 351, y => 237),
  (x => 352, y => 237),
  (x => 353, y => 237),
  (x => 358, y => 237),
  (x => 359, y => 237),
  (x => 360, y => 237),
  (x => 367, y => 237),
  (x => 368, y => 237),
  (x => 369, y => 237),
  (x => 370, y => 237),
  (x => 376, y => 237),
  (x => 377, y => 237),
  (x => 378, y => 237),
  (x => 379, y => 237),
  (x => 386, y => 237),
  (x => 387, y => 237),
  (x => 388, y => 237),
  (x => 389, y => 237),
  (x => 394, y => 237),
  (x => 395, y => 237),
  (x => 396, y => 237),
  (x => 397, y => 237),
  (x => 209, y => 238),
  (x => 210, y => 238),
  (x => 211, y => 238),
  (x => 212, y => 238),
  (x => 213, y => 238),
  (x => 214, y => 238),
  (x => 215, y => 238),
  (x => 216, y => 238),
  (x => 217, y => 238),
  (x => 218, y => 238),
  (x => 219, y => 238),
  (x => 220, y => 238),
  (x => 221, y => 238),
  (x => 228, y => 238),
  (x => 229, y => 238),
  (x => 230, y => 238),
  (x => 231, y => 238),
  (x => 246, y => 238),
  (x => 247, y => 238),
  (x => 248, y => 238),
  (x => 254, y => 238),
  (x => 255, y => 238),
  (x => 256, y => 238),
  (x => 257, y => 238),
  (x => 263, y => 238),
  (x => 264, y => 238),
  (x => 265, y => 238),
  (x => 271, y => 238),
  (x => 272, y => 238),
  (x => 273, y => 238),
  (x => 281, y => 238),
  (x => 282, y => 238),
  (x => 283, y => 238),
  (x => 288, y => 238),
  (x => 289, y => 238),
  (x => 290, y => 238),
  (x => 291, y => 238),
  (x => 317, y => 238),
  (x => 318, y => 238),
  (x => 319, y => 238),
  (x => 320, y => 238),
  (x => 337, y => 238),
  (x => 338, y => 238),
  (x => 339, y => 238),
  (x => 344, y => 238),
  (x => 345, y => 238),
  (x => 346, y => 238),
  (x => 351, y => 238),
  (x => 352, y => 238),
  (x => 353, y => 238),
  (x => 358, y => 238),
  (x => 359, y => 238),
  (x => 367, y => 238),
  (x => 368, y => 238),
  (x => 369, y => 238),
  (x => 370, y => 238),
  (x => 376, y => 238),
  (x => 377, y => 238),
  (x => 378, y => 238),
  (x => 379, y => 238),
  (x => 387, y => 238),
  (x => 388, y => 238),
  (x => 389, y => 238),
  (x => 394, y => 238),
  (x => 395, y => 238),
  (x => 396, y => 238),
  (x => 397, y => 238),
  (x => 209, y => 239),
  (x => 210, y => 239),
  (x => 211, y => 239),
  (x => 212, y => 239),
  (x => 213, y => 239),
  (x => 214, y => 239),
  (x => 215, y => 239),
  (x => 216, y => 239),
  (x => 217, y => 239),
  (x => 218, y => 239),
  (x => 219, y => 239),
  (x => 220, y => 239),
  (x => 221, y => 239),
  (x => 228, y => 239),
  (x => 229, y => 239),
  (x => 230, y => 239),
  (x => 231, y => 239),
  (x => 244, y => 239),
  (x => 245, y => 239),
  (x => 246, y => 239),
  (x => 247, y => 239),
  (x => 248, y => 239),
  (x => 255, y => 239),
  (x => 256, y => 239),
  (x => 257, y => 239),
  (x => 263, y => 239),
  (x => 264, y => 239),
  (x => 270, y => 239),
  (x => 271, y => 239),
  (x => 272, y => 239),
  (x => 273, y => 239),
  (x => 281, y => 239),
  (x => 282, y => 239),
  (x => 283, y => 239),
  (x => 288, y => 239),
  (x => 289, y => 239),
  (x => 290, y => 239),
  (x => 291, y => 239),
  (x => 316, y => 239),
  (x => 317, y => 239),
  (x => 318, y => 239),
  (x => 319, y => 239),
  (x => 337, y => 239),
  (x => 338, y => 239),
  (x => 339, y => 239),
  (x => 340, y => 239),
  (x => 344, y => 239),
  (x => 345, y => 239),
  (x => 346, y => 239),
  (x => 351, y => 239),
  (x => 352, y => 239),
  (x => 353, y => 239),
  (x => 357, y => 239),
  (x => 358, y => 239),
  (x => 359, y => 239),
  (x => 367, y => 239),
  (x => 368, y => 239),
  (x => 369, y => 239),
  (x => 370, y => 239),
  (x => 376, y => 239),
  (x => 377, y => 239),
  (x => 378, y => 239),
  (x => 379, y => 239),
  (x => 387, y => 239),
  (x => 388, y => 239),
  (x => 389, y => 239),
  (x => 395, y => 239),
  (x => 396, y => 239),
  (x => 397, y => 239),
  (x => 398, y => 239),
  (x => 399, y => 239),
  (x => 209, y => 240),
  (x => 210, y => 240),
  (x => 211, y => 240),
  (x => 212, y => 240),
  (x => 213, y => 240),
  (x => 214, y => 240),
  (x => 215, y => 240),
  (x => 216, y => 240),
  (x => 217, y => 240),
  (x => 218, y => 240),
  (x => 219, y => 240),
  (x => 228, y => 240),
  (x => 229, y => 240),
  (x => 230, y => 240),
  (x => 231, y => 240),
  (x => 239, y => 240),
  (x => 240, y => 240),
  (x => 241, y => 240),
  (x => 242, y => 240),
  (x => 243, y => 240),
  (x => 244, y => 240),
  (x => 245, y => 240),
  (x => 246, y => 240),
  (x => 247, y => 240),
  (x => 248, y => 240),
  (x => 255, y => 240),
  (x => 256, y => 240),
  (x => 257, y => 240),
  (x => 262, y => 240),
  (x => 263, y => 240),
  (x => 264, y => 240),
  (x => 270, y => 240),
  (x => 271, y => 240),
  (x => 272, y => 240),
  (x => 273, y => 240),
  (x => 274, y => 240),
  (x => 275, y => 240),
  (x => 276, y => 240),
  (x => 277, y => 240),
  (x => 278, y => 240),
  (x => 279, y => 240),
  (x => 280, y => 240),
  (x => 281, y => 240),
  (x => 282, y => 240),
  (x => 283, y => 240),
  (x => 288, y => 240),
  (x => 289, y => 240),
  (x => 290, y => 240),
  (x => 315, y => 240),
  (x => 316, y => 240),
  (x => 317, y => 240),
  (x => 318, y => 240),
  (x => 338, y => 240),
  (x => 339, y => 240),
  (x => 340, y => 240),
  (x => 344, y => 240),
  (x => 345, y => 240),
  (x => 351, y => 240),
  (x => 352, y => 240),
  (x => 353, y => 240),
  (x => 357, y => 240),
  (x => 358, y => 240),
  (x => 359, y => 240),
  (x => 367, y => 240),
  (x => 368, y => 240),
  (x => 369, y => 240),
  (x => 370, y => 240),
  (x => 376, y => 240),
  (x => 377, y => 240),
  (x => 378, y => 240),
  (x => 379, y => 240),
  (x => 387, y => 240),
  (x => 388, y => 240),
  (x => 389, y => 240),
  (x => 395, y => 240),
  (x => 396, y => 240),
  (x => 397, y => 240),
  (x => 398, y => 240),
  (x => 399, y => 240),
  (x => 400, y => 240),
  (x => 401, y => 240),
  (x => 209, y => 241),
  (x => 210, y => 241),
  (x => 211, y => 241),
  (x => 212, y => 241),
  (x => 213, y => 241),
  (x => 214, y => 241),
  (x => 215, y => 241),
  (x => 216, y => 241),
  (x => 217, y => 241),
  (x => 228, y => 241),
  (x => 229, y => 241),
  (x => 230, y => 241),
  (x => 231, y => 241),
  (x => 238, y => 241),
  (x => 239, y => 241),
  (x => 240, y => 241),
  (x => 241, y => 241),
  (x => 242, y => 241),
  (x => 243, y => 241),
  (x => 244, y => 241),
  (x => 245, y => 241),
  (x => 246, y => 241),
  (x => 247, y => 241),
  (x => 248, y => 241),
  (x => 255, y => 241),
  (x => 256, y => 241),
  (x => 257, y => 241),
  (x => 262, y => 241),
  (x => 263, y => 241),
  (x => 264, y => 241),
  (x => 270, y => 241),
  (x => 271, y => 241),
  (x => 272, y => 241),
  (x => 273, y => 241),
  (x => 274, y => 241),
  (x => 275, y => 241),
  (x => 276, y => 241),
  (x => 277, y => 241),
  (x => 278, y => 241),
  (x => 279, y => 241),
  (x => 280, y => 241),
  (x => 281, y => 241),
  (x => 282, y => 241),
  (x => 283, y => 241),
  (x => 288, y => 241),
  (x => 289, y => 241),
  (x => 290, y => 241),
  (x => 314, y => 241),
  (x => 315, y => 241),
  (x => 316, y => 241),
  (x => 317, y => 241),
  (x => 338, y => 241),
  (x => 339, y => 241),
  (x => 340, y => 241),
  (x => 344, y => 241),
  (x => 345, y => 241),
  (x => 352, y => 241),
  (x => 353, y => 241),
  (x => 354, y => 241),
  (x => 357, y => 241),
  (x => 358, y => 241),
  (x => 359, y => 241),
  (x => 367, y => 241),
  (x => 368, y => 241),
  (x => 369, y => 241),
  (x => 370, y => 241),
  (x => 376, y => 241),
  (x => 377, y => 241),
  (x => 378, y => 241),
  (x => 379, y => 241),
  (x => 387, y => 241),
  (x => 388, y => 241),
  (x => 389, y => 241),
  (x => 396, y => 241),
  (x => 397, y => 241),
  (x => 398, y => 241),
  (x => 399, y => 241),
  (x => 400, y => 241),
  (x => 401, y => 241),
  (x => 402, y => 241),
  (x => 209, y => 242),
  (x => 210, y => 242),
  (x => 211, y => 242),
  (x => 212, y => 242),
  (x => 228, y => 242),
  (x => 229, y => 242),
  (x => 230, y => 242),
  (x => 231, y => 242),
  (x => 237, y => 242),
  (x => 238, y => 242),
  (x => 239, y => 242),
  (x => 240, y => 242),
  (x => 246, y => 242),
  (x => 247, y => 242),
  (x => 248, y => 242),
  (x => 256, y => 242),
  (x => 257, y => 242),
  (x => 258, y => 242),
  (x => 262, y => 242),
  (x => 263, y => 242),
  (x => 264, y => 242),
  (x => 270, y => 242),
  (x => 271, y => 242),
  (x => 272, y => 242),
  (x => 273, y => 242),
  (x => 274, y => 242),
  (x => 275, y => 242),
  (x => 276, y => 242),
  (x => 277, y => 242),
  (x => 278, y => 242),
  (x => 279, y => 242),
  (x => 280, y => 242),
  (x => 281, y => 242),
  (x => 282, y => 242),
  (x => 283, y => 242),
  (x => 288, y => 242),
  (x => 289, y => 242),
  (x => 290, y => 242),
  (x => 313, y => 242),
  (x => 314, y => 242),
  (x => 315, y => 242),
  (x => 316, y => 242),
  (x => 338, y => 242),
  (x => 339, y => 242),
  (x => 340, y => 242),
  (x => 343, y => 242),
  (x => 344, y => 242),
  (x => 345, y => 242),
  (x => 352, y => 242),
  (x => 353, y => 242),
  (x => 354, y => 242),
  (x => 357, y => 242),
  (x => 358, y => 242),
  (x => 359, y => 242),
  (x => 367, y => 242),
  (x => 368, y => 242),
  (x => 369, y => 242),
  (x => 370, y => 242),
  (x => 376, y => 242),
  (x => 377, y => 242),
  (x => 378, y => 242),
  (x => 379, y => 242),
  (x => 387, y => 242),
  (x => 388, y => 242),
  (x => 389, y => 242),
  (x => 397, y => 242),
  (x => 398, y => 242),
  (x => 399, y => 242),
  (x => 400, y => 242),
  (x => 401, y => 242),
  (x => 402, y => 242),
  (x => 403, y => 242),
  (x => 209, y => 243),
  (x => 210, y => 243),
  (x => 211, y => 243),
  (x => 212, y => 243),
  (x => 228, y => 243),
  (x => 229, y => 243),
  (x => 230, y => 243),
  (x => 231, y => 243),
  (x => 237, y => 243),
  (x => 238, y => 243),
  (x => 239, y => 243),
  (x => 246, y => 243),
  (x => 247, y => 243),
  (x => 248, y => 243),
  (x => 256, y => 243),
  (x => 257, y => 243),
  (x => 258, y => 243),
  (x => 262, y => 243),
  (x => 263, y => 243),
  (x => 270, y => 243),
  (x => 271, y => 243),
  (x => 272, y => 243),
  (x => 273, y => 243),
  (x => 288, y => 243),
  (x => 289, y => 243),
  (x => 290, y => 243),
  (x => 312, y => 243),
  (x => 313, y => 243),
  (x => 314, y => 243),
  (x => 315, y => 243),
  (x => 338, y => 243),
  (x => 339, y => 243),
  (x => 340, y => 243),
  (x => 343, y => 243),
  (x => 344, y => 243),
  (x => 345, y => 243),
  (x => 352, y => 243),
  (x => 353, y => 243),
  (x => 354, y => 243),
  (x => 357, y => 243),
  (x => 358, y => 243),
  (x => 367, y => 243),
  (x => 368, y => 243),
  (x => 369, y => 243),
  (x => 370, y => 243),
  (x => 376, y => 243),
  (x => 377, y => 243),
  (x => 378, y => 243),
  (x => 379, y => 243),
  (x => 387, y => 243),
  (x => 388, y => 243),
  (x => 389, y => 243),
  (x => 399, y => 243),
  (x => 400, y => 243),
  (x => 401, y => 243),
  (x => 402, y => 243),
  (x => 403, y => 243),
  (x => 404, y => 243),
  (x => 209, y => 244),
  (x => 210, y => 244),
  (x => 211, y => 244),
  (x => 212, y => 244),
  (x => 228, y => 244),
  (x => 229, y => 244),
  (x => 230, y => 244),
  (x => 231, y => 244),
  (x => 236, y => 244),
  (x => 237, y => 244),
  (x => 238, y => 244),
  (x => 246, y => 244),
  (x => 247, y => 244),
  (x => 248, y => 244),
  (x => 256, y => 244),
  (x => 257, y => 244),
  (x => 258, y => 244),
  (x => 261, y => 244),
  (x => 262, y => 244),
  (x => 263, y => 244),
  (x => 270, y => 244),
  (x => 271, y => 244),
  (x => 272, y => 244),
  (x => 273, y => 244),
  (x => 288, y => 244),
  (x => 289, y => 244),
  (x => 290, y => 244),
  (x => 312, y => 244),
  (x => 313, y => 244),
  (x => 314, y => 244),
  (x => 338, y => 244),
  (x => 339, y => 244),
  (x => 340, y => 244),
  (x => 343, y => 244),
  (x => 344, y => 244),
  (x => 345, y => 244),
  (x => 352, y => 244),
  (x => 353, y => 244),
  (x => 354, y => 244),
  (x => 357, y => 244),
  (x => 358, y => 244),
  (x => 367, y => 244),
  (x => 368, y => 244),
  (x => 369, y => 244),
  (x => 370, y => 244),
  (x => 376, y => 244),
  (x => 377, y => 244),
  (x => 378, y => 244),
  (x => 379, y => 244),
  (x => 387, y => 244),
  (x => 388, y => 244),
  (x => 389, y => 244),
  (x => 401, y => 244),
  (x => 402, y => 244),
  (x => 403, y => 244),
  (x => 404, y => 244),
  (x => 209, y => 245),
  (x => 210, y => 245),
  (x => 211, y => 245),
  (x => 212, y => 245),
  (x => 228, y => 245),
  (x => 229, y => 245),
  (x => 230, y => 245),
  (x => 231, y => 245),
  (x => 236, y => 245),
  (x => 237, y => 245),
  (x => 238, y => 245),
  (x => 246, y => 245),
  (x => 247, y => 245),
  (x => 248, y => 245),
  (x => 257, y => 245),
  (x => 258, y => 245),
  (x => 261, y => 245),
  (x => 262, y => 245),
  (x => 263, y => 245),
  (x => 271, y => 245),
  (x => 272, y => 245),
  (x => 273, y => 245),
  (x => 288, y => 245),
  (x => 289, y => 245),
  (x => 290, y => 245),
  (x => 311, y => 245),
  (x => 312, y => 245),
  (x => 313, y => 245),
  (x => 338, y => 245),
  (x => 339, y => 245),
  (x => 340, y => 245),
  (x => 343, y => 245),
  (x => 344, y => 245),
  (x => 352, y => 245),
  (x => 353, y => 245),
  (x => 354, y => 245),
  (x => 357, y => 245),
  (x => 358, y => 245),
  (x => 367, y => 245),
  (x => 368, y => 245),
  (x => 369, y => 245),
  (x => 370, y => 245),
  (x => 376, y => 245),
  (x => 377, y => 245),
  (x => 378, y => 245),
  (x => 379, y => 245),
  (x => 387, y => 245),
  (x => 388, y => 245),
  (x => 389, y => 245),
  (x => 402, y => 245),
  (x => 403, y => 245),
  (x => 404, y => 245),
  (x => 209, y => 246),
  (x => 210, y => 246),
  (x => 211, y => 246),
  (x => 212, y => 246),
  (x => 228, y => 246),
  (x => 229, y => 246),
  (x => 230, y => 246),
  (x => 231, y => 246),
  (x => 236, y => 246),
  (x => 237, y => 246),
  (x => 238, y => 246),
  (x => 245, y => 246),
  (x => 246, y => 246),
  (x => 247, y => 246),
  (x => 248, y => 246),
  (x => 257, y => 246),
  (x => 258, y => 246),
  (x => 261, y => 246),
  (x => 262, y => 246),
  (x => 271, y => 246),
  (x => 272, y => 246),
  (x => 273, y => 246),
  (x => 288, y => 246),
  (x => 289, y => 246),
  (x => 290, y => 246),
  (x => 311, y => 246),
  (x => 312, y => 246),
  (x => 313, y => 246),
  (x => 339, y => 246),
  (x => 340, y => 246),
  (x => 341, y => 246),
  (x => 342, y => 246),
  (x => 343, y => 246),
  (x => 344, y => 246),
  (x => 353, y => 246),
  (x => 354, y => 246),
  (x => 355, y => 246),
  (x => 356, y => 246),
  (x => 357, y => 246),
  (x => 358, y => 246),
  (x => 367, y => 246),
  (x => 368, y => 246),
  (x => 369, y => 246),
  (x => 370, y => 246),
  (x => 376, y => 246),
  (x => 377, y => 246),
  (x => 378, y => 246),
  (x => 379, y => 246),
  (x => 387, y => 246),
  (x => 388, y => 246),
  (x => 389, y => 246),
  (x => 402, y => 246),
  (x => 403, y => 246),
  (x => 404, y => 246),
  (x => 209, y => 247),
  (x => 210, y => 247),
  (x => 211, y => 247),
  (x => 212, y => 247),
  (x => 228, y => 247),
  (x => 229, y => 247),
  (x => 230, y => 247),
  (x => 231, y => 247),
  (x => 236, y => 247),
  (x => 237, y => 247),
  (x => 238, y => 247),
  (x => 239, y => 247),
  (x => 245, y => 247),
  (x => 246, y => 247),
  (x => 247, y => 247),
  (x => 248, y => 247),
  (x => 257, y => 247),
  (x => 258, y => 247),
  (x => 259, y => 247),
  (x => 260, y => 247),
  (x => 261, y => 247),
  (x => 262, y => 247),
  (x => 271, y => 247),
  (x => 272, y => 247),
  (x => 273, y => 247),
  (x => 274, y => 247),
  (x => 288, y => 247),
  (x => 289, y => 247),
  (x => 290, y => 247),
  (x => 310, y => 247),
  (x => 311, y => 247),
  (x => 312, y => 247),
  (x => 313, y => 247),
  (x => 339, y => 247),
  (x => 340, y => 247),
  (x => 341, y => 247),
  (x => 342, y => 247),
  (x => 343, y => 247),
  (x => 344, y => 247),
  (x => 353, y => 247),
  (x => 354, y => 247),
  (x => 355, y => 247),
  (x => 356, y => 247),
  (x => 357, y => 247),
  (x => 358, y => 247),
  (x => 367, y => 247),
  (x => 368, y => 247),
  (x => 369, y => 247),
  (x => 370, y => 247),
  (x => 376, y => 247),
  (x => 377, y => 247),
  (x => 378, y => 247),
  (x => 379, y => 247),
  (x => 387, y => 247),
  (x => 388, y => 247),
  (x => 389, y => 247),
  (x => 402, y => 247),
  (x => 403, y => 247),
  (x => 404, y => 247),
  (x => 209, y => 248),
  (x => 210, y => 248),
  (x => 211, y => 248),
  (x => 212, y => 248),
  (x => 228, y => 248),
  (x => 229, y => 248),
  (x => 230, y => 248),
  (x => 231, y => 248),
  (x => 236, y => 248),
  (x => 237, y => 248),
  (x => 238, y => 248),
  (x => 239, y => 248),
  (x => 240, y => 248),
  (x => 243, y => 248),
  (x => 244, y => 248),
  (x => 245, y => 248),
  (x => 246, y => 248),
  (x => 247, y => 248),
  (x => 248, y => 248),
  (x => 257, y => 248),
  (x => 258, y => 248),
  (x => 259, y => 248),
  (x => 260, y => 248),
  (x => 261, y => 248),
  (x => 262, y => 248),
  (x => 272, y => 248),
  (x => 273, y => 248),
  (x => 274, y => 248),
  (x => 275, y => 248),
  (x => 276, y => 248),
  (x => 281, y => 248),
  (x => 288, y => 248),
  (x => 289, y => 248),
  (x => 290, y => 248),
  (x => 310, y => 248),
  (x => 311, y => 248),
  (x => 312, y => 248),
  (x => 313, y => 248),
  (x => 339, y => 248),
  (x => 340, y => 248),
  (x => 341, y => 248),
  (x => 342, y => 248),
  (x => 343, y => 248),
  (x => 344, y => 248),
  (x => 353, y => 248),
  (x => 354, y => 248),
  (x => 355, y => 248),
  (x => 356, y => 248),
  (x => 357, y => 248),
  (x => 367, y => 248),
  (x => 368, y => 248),
  (x => 369, y => 248),
  (x => 370, y => 248),
  (x => 376, y => 248),
  (x => 377, y => 248),
  (x => 378, y => 248),
  (x => 379, y => 248),
  (x => 387, y => 248),
  (x => 388, y => 248),
  (x => 389, y => 248),
  (x => 394, y => 248),
  (x => 395, y => 248),
  (x => 401, y => 248),
  (x => 402, y => 248),
  (x => 403, y => 248),
  (x => 404, y => 248),
  (x => 209, y => 249),
  (x => 210, y => 249),
  (x => 211, y => 249),
  (x => 212, y => 249),
  (x => 228, y => 249),
  (x => 229, y => 249),
  (x => 230, y => 249),
  (x => 231, y => 249),
  (x => 237, y => 249),
  (x => 238, y => 249),
  (x => 239, y => 249),
  (x => 240, y => 249),
  (x => 241, y => 249),
  (x => 242, y => 249),
  (x => 243, y => 249),
  (x => 246, y => 249),
  (x => 247, y => 249),
  (x => 248, y => 249),
  (x => 258, y => 249),
  (x => 259, y => 249),
  (x => 260, y => 249),
  (x => 261, y => 249),
  (x => 262, y => 249),
  (x => 272, y => 249),
  (x => 273, y => 249),
  (x => 274, y => 249),
  (x => 275, y => 249),
  (x => 276, y => 249),
  (x => 277, y => 249),
  (x => 278, y => 249),
  (x => 279, y => 249),
  (x => 280, y => 249),
  (x => 281, y => 249),
  (x => 288, y => 249),
  (x => 289, y => 249),
  (x => 290, y => 249),
  (x => 310, y => 249),
  (x => 311, y => 249),
  (x => 312, y => 249),
  (x => 313, y => 249),
  (x => 314, y => 249),
  (x => 315, y => 249),
  (x => 316, y => 249),
  (x => 317, y => 249),
  (x => 318, y => 249),
  (x => 319, y => 249),
  (x => 320, y => 249),
  (x => 321, y => 249),
  (x => 322, y => 249),
  (x => 339, y => 249),
  (x => 340, y => 249),
  (x => 341, y => 249),
  (x => 342, y => 249),
  (x => 343, y => 249),
  (x => 353, y => 249),
  (x => 354, y => 249),
  (x => 355, y => 249),
  (x => 356, y => 249),
  (x => 357, y => 249),
  (x => 367, y => 249),
  (x => 368, y => 249),
  (x => 369, y => 249),
  (x => 370, y => 249),
  (x => 376, y => 249),
  (x => 377, y => 249),
  (x => 378, y => 249),
  (x => 379, y => 249),
  (x => 387, y => 249),
  (x => 388, y => 249),
  (x => 389, y => 249),
  (x => 394, y => 249),
  (x => 395, y => 249),
  (x => 396, y => 249),
  (x => 397, y => 249),
  (x => 398, y => 249),
  (x => 399, y => 249),
  (x => 400, y => 249),
  (x => 401, y => 249),
  (x => 402, y => 249),
  (x => 403, y => 249),
  (x => 209, y => 250),
  (x => 210, y => 250),
  (x => 211, y => 250),
  (x => 212, y => 250),
  (x => 228, y => 250),
  (x => 229, y => 250),
  (x => 230, y => 250),
  (x => 231, y => 250),
  (x => 237, y => 250),
  (x => 238, y => 250),
  (x => 239, y => 250),
  (x => 240, y => 250),
  (x => 241, y => 250),
  (x => 242, y => 250),
  (x => 246, y => 250),
  (x => 247, y => 250),
  (x => 248, y => 250),
  (x => 258, y => 250),
  (x => 259, y => 250),
  (x => 260, y => 250),
  (x => 261, y => 250),
  (x => 273, y => 250),
  (x => 274, y => 250),
  (x => 275, y => 250),
  (x => 276, y => 250),
  (x => 277, y => 250),
  (x => 278, y => 250),
  (x => 279, y => 250),
  (x => 280, y => 250),
  (x => 281, y => 250),
  (x => 288, y => 250),
  (x => 289, y => 250),
  (x => 290, y => 250),
  (x => 310, y => 250),
  (x => 311, y => 250),
  (x => 312, y => 250),
  (x => 313, y => 250),
  (x => 314, y => 250),
  (x => 315, y => 250),
  (x => 316, y => 250),
  (x => 317, y => 250),
  (x => 318, y => 250),
  (x => 319, y => 250),
  (x => 320, y => 250),
  (x => 321, y => 250),
  (x => 322, y => 250),
  (x => 339, y => 250),
  (x => 340, y => 250),
  (x => 341, y => 250),
  (x => 342, y => 250),
  (x => 343, y => 250),
  (x => 353, y => 250),
  (x => 354, y => 250),
  (x => 355, y => 250),
  (x => 356, y => 250),
  (x => 357, y => 250),
  (x => 367, y => 250),
  (x => 368, y => 250),
  (x => 369, y => 250),
  (x => 370, y => 250),
  (x => 376, y => 250),
  (x => 377, y => 250),
  (x => 378, y => 250),
  (x => 379, y => 250),
  (x => 387, y => 250),
  (x => 388, y => 250),
  (x => 389, y => 250),
  (x => 394, y => 250),
  (x => 395, y => 250),
  (x => 396, y => 250),
  (x => 397, y => 250),
  (x => 398, y => 250),
  (x => 399, y => 250),
  (x => 400, y => 250),
  (x => 401, y => 250),
  (x => 402, y => 250),
  (x => 209, y => 251),
  (x => 210, y => 251),
  (x => 211, y => 251),
  (x => 212, y => 251),
  (x => 228, y => 251),
  (x => 229, y => 251),
  (x => 230, y => 251),
  (x => 231, y => 251),
  (x => 238, y => 251),
  (x => 239, y => 251),
  (x => 240, y => 251),
  (x => 241, y => 251),
  (x => 246, y => 251),
  (x => 247, y => 251),
  (x => 248, y => 251),
  (x => 258, y => 251),
  (x => 259, y => 251),
  (x => 260, y => 251),
  (x => 261, y => 251),
  (x => 275, y => 251),
  (x => 276, y => 251),
  (x => 277, y => 251),
  (x => 278, y => 251),
  (x => 279, y => 251),
  (x => 280, y => 251),
  (x => 288, y => 251),
  (x => 289, y => 251),
  (x => 290, y => 251),
  (x => 291, y => 251),
  (x => 310, y => 251),
  (x => 311, y => 251),
  (x => 312, y => 251),
  (x => 313, y => 251),
  (x => 314, y => 251),
  (x => 315, y => 251),
  (x => 316, y => 251),
  (x => 317, y => 251),
  (x => 318, y => 251),
  (x => 319, y => 251),
  (x => 320, y => 251),
  (x => 321, y => 251),
  (x => 322, y => 251),
  (x => 340, y => 251),
  (x => 341, y => 251),
  (x => 342, y => 251),
  (x => 343, y => 251),
  (x => 353, y => 251),
  (x => 354, y => 251),
  (x => 355, y => 251),
  (x => 356, y => 251),
  (x => 357, y => 251),
  (x => 367, y => 251),
  (x => 368, y => 251),
  (x => 369, y => 251),
  (x => 370, y => 251),
  (x => 376, y => 251),
  (x => 377, y => 251),
  (x => 378, y => 251),
  (x => 379, y => 251),
  (x => 387, y => 251),
  (x => 388, y => 251),
  (x => 389, y => 251),
  (x => 395, y => 251),
  (x => 396, y => 251),
  (x => 397, y => 251),
  (x => 398, y => 251),
  (x => 399, y => 251),
  (x => 400, y => 251),
  (x => 401, y => 251),
  (x => 258, y => 252),
  (x => 259, y => 252),
  (x => 260, y => 252),
  (x => 261, y => 252),
  (x => 310, y => 252),
  (x => 311, y => 252),
  (x => 312, y => 252),
  (x => 313, y => 252),
  (x => 314, y => 252),
  (x => 315, y => 252),
  (x => 316, y => 252),
  (x => 317, y => 252),
  (x => 318, y => 252),
  (x => 319, y => 252),
  (x => 320, y => 252),
  (x => 321, y => 252),
  (x => 322, y => 252),
  (x => 258, y => 253),
  (x => 259, y => 253),
  (x => 260, y => 253),
  (x => 258, y => 254),
  (x => 259, y => 254),
  (x => 260, y => 254),
  (x => 258, y => 255),
  (x => 259, y => 255),
  (x => 260, y => 255),
  (x => 257, y => 256),
  (x => 258, y => 256),
  (x => 259, y => 256),
  (x => 256, y => 257),
  (x => 257, y => 257),
  (x => 258, y => 257),
  (x => 259, y => 257),
  (x => 253, y => 258),
  (x => 254, y => 258),
  (x => 255, y => 258),
  (x => 256, y => 258),
  (x => 257, y => 258),
  (x => 258, y => 258),
  (x => 259, y => 258),
  (x => 253, y => 259),
  (x => 254, y => 259),
  (x => 255, y => 259),
  (x => 256, y => 259),
  (x => 257, y => 259),
  (x => 258, y => 259),
  (x => 253, y => 260),
  (x => 254, y => 260),
  (x => 255, y => 260),
  (x => 256, y => 260),
  (x => 257, y => 260),
  (x => 254, y => 261),
  (x => 255, y => 261)
);
	
constant p1_1: CoordPairArray(0 to 112) := (
  (x => 208, y => 26),
  (x => 209, y => 26),
  (x => 210, y => 26),
  (x => 206, y => 27),
  (x => 207, y => 27),
  (x => 208, y => 27),
  (x => 209, y => 27),
  (x => 210, y => 27),
  (x => 204, y => 28),
  (x => 205, y => 28),
  (x => 206, y => 28),
  (x => 207, y => 28),
  (x => 208, y => 28),
  (x => 209, y => 28),
  (x => 210, y => 28),
  (x => 203, y => 29),
  (x => 204, y => 29),
  (x => 205, y => 29),
  (x => 206, y => 29),
  (x => 207, y => 29),
  (x => 208, y => 29),
  (x => 209, y => 29),
  (x => 210, y => 29),
  (x => 203, y => 30),
  (x => 204, y => 30),
  (x => 205, y => 30),
  (x => 206, y => 30),
  (x => 207, y => 30),
  (x => 208, y => 30),
  (x => 209, y => 30),
  (x => 210, y => 30),
  (x => 203, y => 31),
  (x => 204, y => 31),
  (x => 205, y => 31),
  (x => 206, y => 31),
  (x => 207, y => 31),
  (x => 208, y => 31),
  (x => 209, y => 31),
  (x => 210, y => 31),
  (x => 203, y => 32),
  (x => 204, y => 32),
  (x => 207, y => 32),
  (x => 208, y => 32),
  (x => 209, y => 32),
  (x => 210, y => 32),
  (x => 207, y => 33),
  (x => 208, y => 33),
  (x => 209, y => 33),
  (x => 210, y => 33),
  (x => 207, y => 34),
  (x => 208, y => 34),
  (x => 209, y => 34),
  (x => 210, y => 34),
  (x => 207, y => 35),
  (x => 208, y => 35),
  (x => 209, y => 35),
  (x => 210, y => 35),
  (x => 207, y => 36),
  (x => 208, y => 36),
  (x => 209, y => 36),
  (x => 210, y => 36),
  (x => 207, y => 37),
  (x => 208, y => 37),
  (x => 209, y => 37),
  (x => 210, y => 37),
  (x => 207, y => 38),
  (x => 208, y => 38),
  (x => 209, y => 38),
  (x => 210, y => 38),
  (x => 207, y => 39),
  (x => 208, y => 39),
  (x => 209, y => 39),
  (x => 210, y => 39),
  (x => 207, y => 40),
  (x => 208, y => 40),
  (x => 209, y => 40),
  (x => 210, y => 40),
  (x => 207, y => 41),
  (x => 208, y => 41),
  (x => 209, y => 41),
  (x => 210, y => 41),
  (x => 207, y => 42),
  (x => 208, y => 42),
  (x => 209, y => 42),
  (x => 210, y => 42),
  (x => 207, y => 43),
  (x => 208, y => 43),
  (x => 209, y => 43),
  (x => 210, y => 43),
  (x => 207, y => 44),
  (x => 208, y => 44),
  (x => 209, y => 44),
  (x => 210, y => 44),
  (x => 207, y => 45),
  (x => 208, y => 45),
  (x => 209, y => 45),
  (x => 210, y => 45),
  (x => 207, y => 46),
  (x => 208, y => 46),
  (x => 209, y => 46),
  (x => 210, y => 46),
  (x => 207, y => 47),
  (x => 208, y => 47),
  (x => 209, y => 47),
  (x => 210, y => 47),
  (x => 207, y => 48),
  (x => 208, y => 48),
  (x => 209, y => 48),
  (x => 210, y => 48),
  (x => 207, y => 49),
  (x => 208, y => 49),
  (x => 209, y => 49),
  (x => 210, y => 49)
);
constant p1_2: CoordPairArray(0 to 166) := (
  (x => 206, y => 29),
  (x => 207, y => 29),
  (x => 208, y => 29),
  (x => 209, y => 29),
  (x => 210, y => 29),
  (x => 211, y => 29),
  (x => 212, y => 29),
  (x => 205, y => 30),
  (x => 206, y => 30),
  (x => 207, y => 30),
  (x => 208, y => 30),
  (x => 209, y => 30),
  (x => 210, y => 30),
  (x => 211, y => 30),
  (x => 212, y => 30),
  (x => 213, y => 30),
  (x => 205, y => 31),
  (x => 206, y => 31),
  (x => 207, y => 31),
  (x => 208, y => 31),
  (x => 209, y => 31),
  (x => 210, y => 31),
  (x => 211, y => 31),
  (x => 212, y => 31),
  (x => 213, y => 31),
  (x => 214, y => 31),
  (x => 205, y => 32),
  (x => 206, y => 32),
  (x => 207, y => 32),
  (x => 208, y => 32),
  (x => 209, y => 32),
  (x => 210, y => 32),
  (x => 211, y => 32),
  (x => 212, y => 32),
  (x => 213, y => 32),
  (x => 214, y => 32),
  (x => 205, y => 33),
  (x => 206, y => 33),
  (x => 210, y => 33),
  (x => 211, y => 33),
  (x => 212, y => 33),
  (x => 213, y => 33),
  (x => 214, y => 33),
  (x => 211, y => 34),
  (x => 212, y => 34),
  (x => 213, y => 34),
  (x => 214, y => 34),
  (x => 215, y => 34),
  (x => 211, y => 35),
  (x => 212, y => 35),
  (x => 213, y => 35),
  (x => 214, y => 35),
  (x => 215, y => 35),
  (x => 211, y => 36),
  (x => 212, y => 36),
  (x => 213, y => 36),
  (x => 214, y => 36),
  (x => 215, y => 36),
  (x => 211, y => 37),
  (x => 212, y => 37),
  (x => 213, y => 37),
  (x => 214, y => 37),
  (x => 211, y => 38),
  (x => 212, y => 38),
  (x => 213, y => 38),
  (x => 214, y => 38),
  (x => 210, y => 39),
  (x => 211, y => 39),
  (x => 212, y => 39),
  (x => 213, y => 39),
  (x => 214, y => 39),
  (x => 209, y => 40),
  (x => 210, y => 40),
  (x => 211, y => 40),
  (x => 212, y => 40),
  (x => 213, y => 40),
  (x => 208, y => 41),
  (x => 209, y => 41),
  (x => 210, y => 41),
  (x => 211, y => 41),
  (x => 212, y => 41),
  (x => 213, y => 41),
  (x => 207, y => 42),
  (x => 208, y => 42),
  (x => 209, y => 42),
  (x => 210, y => 42),
  (x => 211, y => 42),
  (x => 212, y => 42),
  (x => 207, y => 43),
  (x => 208, y => 43),
  (x => 209, y => 43),
  (x => 210, y => 43),
  (x => 206, y => 44),
  (x => 207, y => 44),
  (x => 208, y => 44),
  (x => 209, y => 44),
  (x => 205, y => 45),
  (x => 206, y => 45),
  (x => 207, y => 45),
  (x => 208, y => 45),
  (x => 205, y => 46),
  (x => 206, y => 46),
  (x => 207, y => 46),
  (x => 204, y => 47),
  (x => 205, y => 47),
  (x => 206, y => 47),
  (x => 207, y => 47),
  (x => 204, y => 48),
  (x => 205, y => 48),
  (x => 206, y => 48),
  (x => 207, y => 48),
  (x => 208, y => 48),
  (x => 209, y => 48),
  (x => 210, y => 48),
  (x => 211, y => 48),
  (x => 212, y => 48),
  (x => 213, y => 48),
  (x => 214, y => 48),
  (x => 215, y => 48),
  (x => 204, y => 49),
  (x => 205, y => 49),
  (x => 206, y => 49),
  (x => 207, y => 49),
  (x => 208, y => 49),
  (x => 209, y => 49),
  (x => 210, y => 49),
  (x => 211, y => 49),
  (x => 212, y => 49),
  (x => 213, y => 49),
  (x => 214, y => 49),
  (x => 215, y => 49),
  (x => 204, y => 50),
  (x => 205, y => 50),
  (x => 206, y => 50),
  (x => 207, y => 50),
  (x => 208, y => 50),
  (x => 209, y => 50),
  (x => 210, y => 50),
  (x => 211, y => 50),
  (x => 212, y => 50),
  (x => 213, y => 50),
  (x => 214, y => 50),
  (x => 215, y => 50),
  (x => 204, y => 51),
  (x => 205, y => 51),
  (x => 206, y => 51),
  (x => 207, y => 51),
  (x => 208, y => 51),
  (x => 209, y => 51),
  (x => 210, y => 51),
  (x => 211, y => 51),
  (x => 212, y => 51),
  (x => 213, y => 51),
  (x => 214, y => 51),
  (x => 215, y => 51),
  (x => 204, y => 52),
  (x => 205, y => 52),
  (x => 206, y => 52),
  (x => 207, y => 52),
  (x => 208, y => 52),
  (x => 209, y => 52),
  (x => 210, y => 52),
  (x => 211, y => 52),
  (x => 212, y => 52),
  (x => 213, y => 52),
  (x => 214, y => 52),
  (x => 215, y => 52)
);
constant p1_3: CoordPairArray(0 to 157) := (
  (x => 204, y => 29),
  (x => 205, y => 29),
  (x => 206, y => 29),
  (x => 207, y => 29),
  (x => 208, y => 29),
  (x => 209, y => 29),
  (x => 210, y => 29),
  (x => 211, y => 29),
  (x => 204, y => 30),
  (x => 205, y => 30),
  (x => 206, y => 30),
  (x => 207, y => 30),
  (x => 208, y => 30),
  (x => 209, y => 30),
  (x => 210, y => 30),
  (x => 211, y => 30),
  (x => 212, y => 30),
  (x => 204, y => 31),
  (x => 205, y => 31),
  (x => 206, y => 31),
  (x => 207, y => 31),
  (x => 208, y => 31),
  (x => 209, y => 31),
  (x => 210, y => 31),
  (x => 211, y => 31),
  (x => 212, y => 31),
  (x => 213, y => 31),
  (x => 204, y => 32),
  (x => 205, y => 32),
  (x => 206, y => 32),
  (x => 207, y => 32),
  (x => 208, y => 32),
  (x => 209, y => 32),
  (x => 210, y => 32),
  (x => 211, y => 32),
  (x => 212, y => 32),
  (x => 213, y => 32),
  (x => 210, y => 33),
  (x => 211, y => 33),
  (x => 212, y => 33),
  (x => 213, y => 33),
  (x => 210, y => 34),
  (x => 211, y => 34),
  (x => 212, y => 34),
  (x => 213, y => 34),
  (x => 210, y => 35),
  (x => 211, y => 35),
  (x => 212, y => 35),
  (x => 213, y => 35),
  (x => 210, y => 36),
  (x => 211, y => 36),
  (x => 212, y => 36),
  (x => 213, y => 36),
  (x => 209, y => 37),
  (x => 210, y => 37),
  (x => 211, y => 37),
  (x => 212, y => 37),
  (x => 213, y => 37),
  (x => 207, y => 38),
  (x => 208, y => 38),
  (x => 209, y => 38),
  (x => 210, y => 38),
  (x => 211, y => 38),
  (x => 212, y => 38),
  (x => 205, y => 39),
  (x => 206, y => 39),
  (x => 207, y => 39),
  (x => 208, y => 39),
  (x => 209, y => 39),
  (x => 210, y => 39),
  (x => 205, y => 40),
  (x => 206, y => 40),
  (x => 207, y => 40),
  (x => 208, y => 40),
  (x => 209, y => 40),
  (x => 210, y => 40),
  (x => 205, y => 41),
  (x => 206, y => 41),
  (x => 207, y => 41),
  (x => 208, y => 41),
  (x => 209, y => 41),
  (x => 210, y => 41),
  (x => 211, y => 41),
  (x => 205, y => 42),
  (x => 206, y => 42),
  (x => 207, y => 42),
  (x => 208, y => 42),
  (x => 209, y => 42),
  (x => 210, y => 42),
  (x => 211, y => 42),
  (x => 212, y => 42),
  (x => 213, y => 42),
  (x => 210, y => 43),
  (x => 211, y => 43),
  (x => 212, y => 43),
  (x => 213, y => 43),
  (x => 210, y => 44),
  (x => 211, y => 44),
  (x => 212, y => 44),
  (x => 213, y => 44),
  (x => 214, y => 44),
  (x => 211, y => 45),
  (x => 212, y => 45),
  (x => 213, y => 45),
  (x => 214, y => 45),
  (x => 211, y => 46),
  (x => 212, y => 46),
  (x => 213, y => 46),
  (x => 214, y => 46),
  (x => 210, y => 47),
  (x => 211, y => 47),
  (x => 212, y => 47),
  (x => 213, y => 47),
  (x => 214, y => 47),
  (x => 203, y => 48),
  (x => 204, y => 48),
  (x => 209, y => 48),
  (x => 210, y => 48),
  (x => 211, y => 48),
  (x => 212, y => 48),
  (x => 213, y => 48),
  (x => 204, y => 49),
  (x => 205, y => 49),
  (x => 206, y => 49),
  (x => 207, y => 49),
  (x => 208, y => 49),
  (x => 209, y => 49),
  (x => 210, y => 49),
  (x => 211, y => 49),
  (x => 212, y => 49),
  (x => 213, y => 49),
  (x => 204, y => 50),
  (x => 205, y => 50),
  (x => 206, y => 50),
  (x => 207, y => 50),
  (x => 208, y => 50),
  (x => 209, y => 50),
  (x => 210, y => 50),
  (x => 211, y => 50),
  (x => 212, y => 50),
  (x => 213, y => 50),
  (x => 203, y => 51),
  (x => 204, y => 51),
  (x => 205, y => 51),
  (x => 206, y => 51),
  (x => 207, y => 51),
  (x => 208, y => 51),
  (x => 209, y => 51),
  (x => 210, y => 51),
  (x => 211, y => 51),
  (x => 212, y => 51),
  (x => 204, y => 52),
  (x => 205, y => 52),
  (x => 206, y => 52),
  (x => 207, y => 52),
  (x => 208, y => 52),
  (x => 209, y => 52),
  (x => 210, y => 52)
);
constant p1_4: CoordPairArray(0 to 150) := (
  (x => 207, y => 31),
  (x => 208, y => 31),
  (x => 209, y => 31),
  (x => 210, y => 31),
  (x => 206, y => 32),
  (x => 207, y => 32),
  (x => 208, y => 32),
  (x => 209, y => 32),
  (x => 210, y => 32),
  (x => 206, y => 33),
  (x => 207, y => 33),
  (x => 208, y => 33),
  (x => 209, y => 33),
  (x => 210, y => 33),
  (x => 206, y => 34),
  (x => 207, y => 34),
  (x => 208, y => 34),
  (x => 209, y => 34),
  (x => 210, y => 34),
  (x => 205, y => 35),
  (x => 206, y => 35),
  (x => 207, y => 35),
  (x => 208, y => 35),
  (x => 209, y => 35),
  (x => 210, y => 35),
  (x => 205, y => 36),
  (x => 206, y => 36),
  (x => 207, y => 36),
  (x => 208, y => 36),
  (x => 209, y => 36),
  (x => 210, y => 36),
  (x => 204, y => 37),
  (x => 205, y => 37),
  (x => 206, y => 37),
  (x => 207, y => 37),
  (x => 208, y => 37),
  (x => 209, y => 37),
  (x => 210, y => 37),
  (x => 204, y => 38),
  (x => 205, y => 38),
  (x => 208, y => 38),
  (x => 209, y => 38),
  (x => 210, y => 38),
  (x => 203, y => 39),
  (x => 204, y => 39),
  (x => 205, y => 39),
  (x => 208, y => 39),
  (x => 209, y => 39),
  (x => 210, y => 39),
  (x => 203, y => 40),
  (x => 204, y => 40),
  (x => 208, y => 40),
  (x => 209, y => 40),
  (x => 210, y => 40),
  (x => 202, y => 41),
  (x => 203, y => 41),
  (x => 204, y => 41),
  (x => 208, y => 41),
  (x => 209, y => 41),
  (x => 210, y => 41),
  (x => 202, y => 42),
  (x => 203, y => 42),
  (x => 208, y => 42),
  (x => 209, y => 42),
  (x => 210, y => 42),
  (x => 201, y => 43),
  (x => 202, y => 43),
  (x => 203, y => 43),
  (x => 208, y => 43),
  (x => 209, y => 43),
  (x => 210, y => 43),
  (x => 200, y => 44),
  (x => 201, y => 44),
  (x => 202, y => 44),
  (x => 208, y => 44),
  (x => 209, y => 44),
  (x => 210, y => 44),
  (x => 200, y => 45),
  (x => 201, y => 45),
  (x => 202, y => 45),
  (x => 208, y => 45),
  (x => 209, y => 45),
  (x => 210, y => 45),
  (x => 200, y => 46),
  (x => 201, y => 46),
  (x => 202, y => 46),
  (x => 204, y => 46),
  (x => 205, y => 46),
  (x => 206, y => 46),
  (x => 207, y => 46),
  (x => 208, y => 46),
  (x => 209, y => 46),
  (x => 210, y => 46),
  (x => 211, y => 46),
  (x => 212, y => 46),
  (x => 213, y => 46),
  (x => 200, y => 47),
  (x => 201, y => 47),
  (x => 202, y => 47),
  (x => 203, y => 47),
  (x => 204, y => 47),
  (x => 205, y => 47),
  (x => 206, y => 47),
  (x => 207, y => 47),
  (x => 208, y => 47),
  (x => 209, y => 47),
  (x => 210, y => 47),
  (x => 211, y => 47),
  (x => 212, y => 47),
  (x => 213, y => 47),
  (x => 200, y => 48),
  (x => 201, y => 48),
  (x => 202, y => 48),
  (x => 203, y => 48),
  (x => 204, y => 48),
  (x => 205, y => 48),
  (x => 206, y => 48),
  (x => 207, y => 48),
  (x => 208, y => 48),
  (x => 209, y => 48),
  (x => 210, y => 48),
  (x => 211, y => 48),
  (x => 212, y => 48),
  (x => 213, y => 48),
  (x => 199, y => 49),
  (x => 200, y => 49),
  (x => 201, y => 49),
  (x => 202, y => 49),
  (x => 203, y => 49),
  (x => 204, y => 49),
  (x => 205, y => 49),
  (x => 206, y => 49),
  (x => 207, y => 49),
  (x => 208, y => 49),
  (x => 209, y => 49),
  (x => 210, y => 49),
  (x => 211, y => 49),
  (x => 212, y => 49),
  (x => 213, y => 49),
  (x => 208, y => 50),
  (x => 209, y => 50),
  (x => 210, y => 50),
  (x => 208, y => 51),
  (x => 209, y => 51),
  (x => 210, y => 51),
  (x => 208, y => 52),
  (x => 209, y => 52),
  (x => 210, y => 52),
  (x => 208, y => 53),
  (x => 209, y => 53),
  (x => 210, y => 53)
);
constant p1_5: CoordPairArray(0 to 167) := (
  (x => 202, y => 29),
  (x => 203, y => 29),
  (x => 204, y => 29),
  (x => 205, y => 29),
  (x => 206, y => 29),
  (x => 207, y => 29),
  (x => 208, y => 29),
  (x => 209, y => 29),
  (x => 210, y => 29),
  (x => 211, y => 29),
  (x => 202, y => 30),
  (x => 203, y => 30),
  (x => 204, y => 30),
  (x => 205, y => 30),
  (x => 206, y => 30),
  (x => 207, y => 30),
  (x => 208, y => 30),
  (x => 209, y => 30),
  (x => 210, y => 30),
  (x => 202, y => 31),
  (x => 203, y => 31),
  (x => 204, y => 31),
  (x => 205, y => 31),
  (x => 206, y => 31),
  (x => 207, y => 31),
  (x => 208, y => 31),
  (x => 209, y => 31),
  (x => 210, y => 31),
  (x => 202, y => 32),
  (x => 203, y => 32),
  (x => 204, y => 32),
  (x => 205, y => 32),
  (x => 206, y => 32),
  (x => 207, y => 32),
  (x => 208, y => 32),
  (x => 209, y => 32),
  (x => 210, y => 32),
  (x => 202, y => 33),
  (x => 203, y => 33),
  (x => 204, y => 33),
  (x => 205, y => 33),
  (x => 206, y => 33),
  (x => 207, y => 33),
  (x => 208, y => 33),
  (x => 209, y => 33),
  (x => 210, y => 33),
  (x => 211, y => 33),
  (x => 202, y => 34),
  (x => 203, y => 34),
  (x => 204, y => 34),
  (x => 202, y => 35),
  (x => 203, y => 35),
  (x => 204, y => 35),
  (x => 202, y => 36),
  (x => 203, y => 36),
  (x => 204, y => 36),
  (x => 202, y => 37),
  (x => 203, y => 37),
  (x => 204, y => 37),
  (x => 202, y => 38),
  (x => 203, y => 38),
  (x => 204, y => 38),
  (x => 205, y => 38),
  (x => 206, y => 38),
  (x => 207, y => 38),
  (x => 208, y => 38),
  (x => 202, y => 39),
  (x => 203, y => 39),
  (x => 204, y => 39),
  (x => 205, y => 39),
  (x => 206, y => 39),
  (x => 207, y => 39),
  (x => 208, y => 39),
  (x => 209, y => 39),
  (x => 210, y => 39),
  (x => 202, y => 40),
  (x => 203, y => 40),
  (x => 204, y => 40),
  (x => 205, y => 40),
  (x => 206, y => 40),
  (x => 207, y => 40),
  (x => 208, y => 40),
  (x => 209, y => 40),
  (x => 210, y => 40),
  (x => 202, y => 41),
  (x => 203, y => 41),
  (x => 204, y => 41),
  (x => 205, y => 41),
  (x => 206, y => 41),
  (x => 207, y => 41),
  (x => 208, y => 41),
  (x => 209, y => 41),
  (x => 210, y => 41),
  (x => 211, y => 41),
  (x => 201, y => 42),
  (x => 202, y => 42),
  (x => 203, y => 42),
  (x => 204, y => 42),
  (x => 205, y => 42),
  (x => 206, y => 42),
  (x => 207, y => 42),
  (x => 208, y => 42),
  (x => 209, y => 42),
  (x => 210, y => 42),
  (x => 211, y => 42),
  (x => 207, y => 43),
  (x => 208, y => 43),
  (x => 209, y => 43),
  (x => 210, y => 43),
  (x => 211, y => 43),
  (x => 208, y => 44),
  (x => 209, y => 44),
  (x => 210, y => 44),
  (x => 211, y => 44),
  (x => 208, y => 45),
  (x => 209, y => 45),
  (x => 210, y => 45),
  (x => 211, y => 45),
  (x => 208, y => 46),
  (x => 209, y => 46),
  (x => 210, y => 46),
  (x => 211, y => 46),
  (x => 208, y => 47),
  (x => 209, y => 47),
  (x => 210, y => 47),
  (x => 211, y => 47),
  (x => 201, y => 48),
  (x => 207, y => 48),
  (x => 208, y => 48),
  (x => 209, y => 48),
  (x => 210, y => 48),
  (x => 211, y => 48),
  (x => 201, y => 49),
  (x => 202, y => 49),
  (x => 203, y => 49),
  (x => 204, y => 49),
  (x => 205, y => 49),
  (x => 206, y => 49),
  (x => 207, y => 49),
  (x => 208, y => 49),
  (x => 209, y => 49),
  (x => 210, y => 49),
  (x => 201, y => 50),
  (x => 202, y => 50),
  (x => 203, y => 50),
  (x => 204, y => 50),
  (x => 205, y => 50),
  (x => 206, y => 50),
  (x => 207, y => 50),
  (x => 208, y => 50),
  (x => 209, y => 50),
  (x => 210, y => 50),
  (x => 201, y => 51),
  (x => 202, y => 51),
  (x => 203, y => 51),
  (x => 204, y => 51),
  (x => 205, y => 51),
  (x => 206, y => 51),
  (x => 207, y => 51),
  (x => 208, y => 51),
  (x => 209, y => 51),
  (x => 201, y => 52),
  (x => 202, y => 52),
  (x => 203, y => 52),
  (x => 204, y => 52),
  (x => 205, y => 52),
  (x => 206, y => 52),
  (x => 207, y => 52)
);
constant p1_6: CoordPairArray(0 to 188) := (
  (x => 208, y => 27),
  (x => 209, y => 27),
  (x => 210, y => 27),
  (x => 211, y => 27),
  (x => 206, y => 28),
  (x => 207, y => 28),
  (x => 208, y => 28),
  (x => 209, y => 28),
  (x => 210, y => 28),
  (x => 211, y => 28),
  (x => 212, y => 28),
  (x => 204, y => 29),
  (x => 205, y => 29),
  (x => 206, y => 29),
  (x => 207, y => 29),
  (x => 208, y => 29),
  (x => 209, y => 29),
  (x => 210, y => 29),
  (x => 211, y => 29),
  (x => 212, y => 29),
  (x => 204, y => 30),
  (x => 205, y => 30),
  (x => 206, y => 30),
  (x => 207, y => 30),
  (x => 208, y => 30),
  (x => 209, y => 30),
  (x => 210, y => 30),
  (x => 211, y => 30),
  (x => 212, y => 30),
  (x => 203, y => 31),
  (x => 204, y => 31),
  (x => 205, y => 31),
  (x => 206, y => 31),
  (x => 207, y => 31),
  (x => 208, y => 31),
  (x => 203, y => 32),
  (x => 204, y => 32),
  (x => 205, y => 32),
  (x => 206, y => 32),
  (x => 202, y => 33),
  (x => 203, y => 33),
  (x => 204, y => 33),
  (x => 205, y => 33),
  (x => 202, y => 34),
  (x => 203, y => 34),
  (x => 204, y => 34),
  (x => 205, y => 34),
  (x => 202, y => 35),
  (x => 203, y => 35),
  (x => 204, y => 35),
  (x => 202, y => 36),
  (x => 203, y => 36),
  (x => 204, y => 36),
  (x => 208, y => 36),
  (x => 209, y => 36),
  (x => 210, y => 36),
  (x => 201, y => 37),
  (x => 202, y => 37),
  (x => 203, y => 37),
  (x => 204, y => 37),
  (x => 207, y => 37),
  (x => 208, y => 37),
  (x => 209, y => 37),
  (x => 210, y => 37),
  (x => 211, y => 37),
  (x => 212, y => 37),
  (x => 201, y => 38),
  (x => 202, y => 38),
  (x => 203, y => 38),
  (x => 204, y => 38),
  (x => 205, y => 38),
  (x => 206, y => 38),
  (x => 207, y => 38),
  (x => 208, y => 38),
  (x => 209, y => 38),
  (x => 210, y => 38),
  (x => 211, y => 38),
  (x => 212, y => 38),
  (x => 201, y => 39),
  (x => 202, y => 39),
  (x => 203, y => 39),
  (x => 204, y => 39),
  (x => 205, y => 39),
  (x => 206, y => 39),
  (x => 207, y => 39),
  (x => 208, y => 39),
  (x => 209, y => 39),
  (x => 210, y => 39),
  (x => 211, y => 39),
  (x => 212, y => 39),
  (x => 201, y => 40),
  (x => 202, y => 40),
  (x => 203, y => 40),
  (x => 204, y => 40),
  (x => 205, y => 40),
  (x => 206, y => 40),
  (x => 209, y => 40),
  (x => 210, y => 40),
  (x => 211, y => 40),
  (x => 212, y => 40),
  (x => 213, y => 40),
  (x => 201, y => 41),
  (x => 202, y => 41),
  (x => 203, y => 41),
  (x => 204, y => 41),
  (x => 205, y => 41),
  (x => 210, y => 41),
  (x => 211, y => 41),
  (x => 212, y => 41),
  (x => 213, y => 41),
  (x => 201, y => 42),
  (x => 202, y => 42),
  (x => 203, y => 42),
  (x => 204, y => 42),
  (x => 205, y => 42),
  (x => 210, y => 42),
  (x => 211, y => 42),
  (x => 212, y => 42),
  (x => 213, y => 42),
  (x => 201, y => 43),
  (x => 202, y => 43),
  (x => 203, y => 43),
  (x => 204, y => 43),
  (x => 210, y => 43),
  (x => 211, y => 43),
  (x => 212, y => 43),
  (x => 213, y => 43),
  (x => 202, y => 44),
  (x => 203, y => 44),
  (x => 204, y => 44),
  (x => 210, y => 44),
  (x => 211, y => 44),
  (x => 212, y => 44),
  (x => 213, y => 44),
  (x => 202, y => 45),
  (x => 203, y => 45),
  (x => 204, y => 45),
  (x => 205, y => 45),
  (x => 210, y => 45),
  (x => 211, y => 45),
  (x => 212, y => 45),
  (x => 213, y => 45),
  (x => 202, y => 46),
  (x => 203, y => 46),
  (x => 204, y => 46),
  (x => 205, y => 46),
  (x => 210, y => 46),
  (x => 211, y => 46),
  (x => 212, y => 46),
  (x => 213, y => 46),
  (x => 202, y => 47),
  (x => 203, y => 47),
  (x => 204, y => 47),
  (x => 205, y => 47),
  (x => 206, y => 47),
  (x => 207, y => 47),
  (x => 208, y => 47),
  (x => 209, y => 47),
  (x => 210, y => 47),
  (x => 211, y => 47),
  (x => 212, y => 47),
  (x => 203, y => 48),
  (x => 204, y => 48),
  (x => 205, y => 48),
  (x => 206, y => 48),
  (x => 207, y => 48),
  (x => 208, y => 48),
  (x => 209, y => 48),
  (x => 210, y => 48),
  (x => 211, y => 48),
  (x => 212, y => 48),
  (x => 203, y => 49),
  (x => 204, y => 49),
  (x => 205, y => 49),
  (x => 206, y => 49),
  (x => 207, y => 49),
  (x => 208, y => 49),
  (x => 209, y => 49),
  (x => 210, y => 49),
  (x => 211, y => 49),
  (x => 204, y => 50),
  (x => 205, y => 50),
  (x => 206, y => 50),
  (x => 207, y => 50),
  (x => 208, y => 50),
  (x => 209, y => 50),
  (x => 210, y => 50),
  (x => 207, y => 51),
  (x => 208, y => 51)
);
constant p1_7: CoordPairArray(0 to 137) := (
  (x => 200, y => 27),
  (x => 201, y => 27),
  (x => 202, y => 27),
  (x => 203, y => 27),
  (x => 204, y => 27),
  (x => 205, y => 27),
  (x => 206, y => 27),
  (x => 207, y => 27),
  (x => 208, y => 27),
  (x => 209, y => 27),
  (x => 210, y => 27),
  (x => 211, y => 27),
  (x => 212, y => 27),
  (x => 200, y => 28),
  (x => 201, y => 28),
  (x => 202, y => 28),
  (x => 203, y => 28),
  (x => 204, y => 28),
  (x => 205, y => 28),
  (x => 206, y => 28),
  (x => 207, y => 28),
  (x => 208, y => 28),
  (x => 209, y => 28),
  (x => 210, y => 28),
  (x => 211, y => 28),
  (x => 212, y => 28),
  (x => 200, y => 29),
  (x => 201, y => 29),
  (x => 202, y => 29),
  (x => 203, y => 29),
  (x => 204, y => 29),
  (x => 205, y => 29),
  (x => 206, y => 29),
  (x => 207, y => 29),
  (x => 208, y => 29),
  (x => 209, y => 29),
  (x => 210, y => 29),
  (x => 211, y => 29),
  (x => 212, y => 29),
  (x => 200, y => 30),
  (x => 201, y => 30),
  (x => 202, y => 30),
  (x => 203, y => 30),
  (x => 204, y => 30),
  (x => 205, y => 30),
  (x => 206, y => 30),
  (x => 207, y => 30),
  (x => 208, y => 30),
  (x => 209, y => 30),
  (x => 210, y => 30),
  (x => 211, y => 30),
  (x => 212, y => 30),
  (x => 200, y => 31),
  (x => 201, y => 31),
  (x => 202, y => 31),
  (x => 203, y => 31),
  (x => 204, y => 31),
  (x => 205, y => 31),
  (x => 206, y => 31),
  (x => 207, y => 31),
  (x => 208, y => 31),
  (x => 209, y => 31),
  (x => 210, y => 31),
  (x => 211, y => 31),
  (x => 208, y => 32),
  (x => 209, y => 32),
  (x => 210, y => 32),
  (x => 211, y => 32),
  (x => 208, y => 33),
  (x => 209, y => 33),
  (x => 210, y => 33),
  (x => 208, y => 34),
  (x => 209, y => 34),
  (x => 210, y => 34),
  (x => 207, y => 35),
  (x => 208, y => 35),
  (x => 209, y => 35),
  (x => 210, y => 35),
  (x => 207, y => 36),
  (x => 208, y => 36),
  (x => 209, y => 36),
  (x => 206, y => 37),
  (x => 207, y => 37),
  (x => 208, y => 37),
  (x => 209, y => 37),
  (x => 206, y => 38),
  (x => 207, y => 38),
  (x => 208, y => 38),
  (x => 209, y => 38),
  (x => 205, y => 39),
  (x => 206, y => 39),
  (x => 207, y => 39),
  (x => 208, y => 39),
  (x => 205, y => 40),
  (x => 206, y => 40),
  (x => 207, y => 40),
  (x => 208, y => 40),
  (x => 205, y => 41),
  (x => 206, y => 41),
  (x => 207, y => 41),
  (x => 208, y => 41),
  (x => 204, y => 42),
  (x => 205, y => 42),
  (x => 206, y => 42),
  (x => 207, y => 42),
  (x => 204, y => 43),
  (x => 205, y => 43),
  (x => 206, y => 43),
  (x => 207, y => 43),
  (x => 204, y => 44),
  (x => 205, y => 44),
  (x => 206, y => 44),
  (x => 207, y => 44),
  (x => 204, y => 45),
  (x => 205, y => 45),
  (x => 206, y => 45),
  (x => 207, y => 45),
  (x => 203, y => 46),
  (x => 204, y => 46),
  (x => 205, y => 46),
  (x => 206, y => 46),
  (x => 207, y => 46),
  (x => 203, y => 47),
  (x => 204, y => 47),
  (x => 205, y => 47),
  (x => 206, y => 47),
  (x => 203, y => 48),
  (x => 204, y => 48),
  (x => 205, y => 48),
  (x => 206, y => 48),
  (x => 203, y => 49),
  (x => 204, y => 49),
  (x => 205, y => 49),
  (x => 206, y => 49),
  (x => 203, y => 50),
  (x => 204, y => 50),
  (x => 205, y => 50),
  (x => 206, y => 50)
);
constant p1_8: CoordPairArray(0 to 191) := (
  (x => 203, y => 23),
  (x => 204, y => 23),
  (x => 205, y => 23),
  (x => 206, y => 23),
  (x => 207, y => 23),
  (x => 208, y => 23),
  (x => 209, y => 23),
  (x => 202, y => 24),
  (x => 203, y => 24),
  (x => 204, y => 24),
  (x => 205, y => 24),
  (x => 206, y => 24),
  (x => 207, y => 24),
  (x => 208, y => 24),
  (x => 209, y => 24),
  (x => 210, y => 24),
  (x => 202, y => 25),
  (x => 203, y => 25),
  (x => 204, y => 25),
  (x => 205, y => 25),
  (x => 206, y => 25),
  (x => 207, y => 25),
  (x => 208, y => 25),
  (x => 209, y => 25),
  (x => 210, y => 25),
  (x => 211, y => 25),
  (x => 201, y => 26),
  (x => 202, y => 26),
  (x => 203, y => 26),
  (x => 204, y => 26),
  (x => 205, y => 26),
  (x => 208, y => 26),
  (x => 209, y => 26),
  (x => 210, y => 26),
  (x => 211, y => 26),
  (x => 201, y => 27),
  (x => 202, y => 27),
  (x => 203, y => 27),
  (x => 204, y => 27),
  (x => 209, y => 27),
  (x => 210, y => 27),
  (x => 211, y => 27),
  (x => 212, y => 27),
  (x => 201, y => 28),
  (x => 202, y => 28),
  (x => 203, y => 28),
  (x => 209, y => 28),
  (x => 210, y => 28),
  (x => 211, y => 28),
  (x => 212, y => 28),
  (x => 201, y => 29),
  (x => 202, y => 29),
  (x => 203, y => 29),
  (x => 209, y => 29),
  (x => 210, y => 29),
  (x => 211, y => 29),
  (x => 212, y => 29),
  (x => 201, y => 30),
  (x => 202, y => 30),
  (x => 203, y => 30),
  (x => 209, y => 30),
  (x => 210, y => 30),
  (x => 211, y => 30),
  (x => 201, y => 31),
  (x => 202, y => 31),
  (x => 203, y => 31),
  (x => 204, y => 31),
  (x => 209, y => 31),
  (x => 210, y => 31),
  (x => 211, y => 31),
  (x => 202, y => 32),
  (x => 203, y => 32),
  (x => 204, y => 32),
  (x => 205, y => 32),
  (x => 207, y => 32),
  (x => 208, y => 32),
  (x => 209, y => 32),
  (x => 210, y => 32),
  (x => 203, y => 33),
  (x => 204, y => 33),
  (x => 205, y => 33),
  (x => 206, y => 33),
  (x => 207, y => 33),
  (x => 208, y => 33),
  (x => 209, y => 33),
  (x => 203, y => 34),
  (x => 204, y => 34),
  (x => 205, y => 34),
  (x => 206, y => 34),
  (x => 207, y => 34),
  (x => 208, y => 34),
  (x => 209, y => 34),
  (x => 203, y => 35),
  (x => 204, y => 35),
  (x => 205, y => 35),
  (x => 206, y => 35),
  (x => 207, y => 35),
  (x => 208, y => 35),
  (x => 209, y => 35),
  (x => 202, y => 36),
  (x => 203, y => 36),
  (x => 204, y => 36),
  (x => 205, y => 36),
  (x => 206, y => 36),
  (x => 207, y => 36),
  (x => 208, y => 36),
  (x => 209, y => 36),
  (x => 210, y => 36),
  (x => 211, y => 36),
  (x => 201, y => 37),
  (x => 202, y => 37),
  (x => 203, y => 37),
  (x => 204, y => 37),
  (x => 209, y => 37),
  (x => 210, y => 37),
  (x => 211, y => 37),
  (x => 201, y => 38),
  (x => 202, y => 38),
  (x => 203, y => 38),
  (x => 209, y => 38),
  (x => 210, y => 38),
  (x => 211, y => 38),
  (x => 212, y => 38),
  (x => 200, y => 39),
  (x => 201, y => 39),
  (x => 202, y => 39),
  (x => 203, y => 39),
  (x => 209, y => 39),
  (x => 210, y => 39),
  (x => 211, y => 39),
  (x => 212, y => 39),
  (x => 200, y => 40),
  (x => 201, y => 40),
  (x => 202, y => 40),
  (x => 203, y => 40),
  (x => 209, y => 40),
  (x => 210, y => 40),
  (x => 211, y => 40),
  (x => 212, y => 40),
  (x => 200, y => 41),
  (x => 201, y => 41),
  (x => 202, y => 41),
  (x => 203, y => 41),
  (x => 209, y => 41),
  (x => 210, y => 41),
  (x => 211, y => 41),
  (x => 212, y => 41),
  (x => 200, y => 42),
  (x => 201, y => 42),
  (x => 202, y => 42),
  (x => 203, y => 42),
  (x => 209, y => 42),
  (x => 210, y => 42),
  (x => 211, y => 42),
  (x => 212, y => 42),
  (x => 201, y => 43),
  (x => 202, y => 43),
  (x => 203, y => 43),
  (x => 204, y => 43),
  (x => 205, y => 43),
  (x => 207, y => 43),
  (x => 208, y => 43),
  (x => 209, y => 43),
  (x => 210, y => 43),
  (x => 211, y => 43),
  (x => 212, y => 43),
  (x => 201, y => 44),
  (x => 202, y => 44),
  (x => 203, y => 44),
  (x => 204, y => 44),
  (x => 205, y => 44),
  (x => 206, y => 44),
  (x => 207, y => 44),
  (x => 208, y => 44),
  (x => 209, y => 44),
  (x => 210, y => 44),
  (x => 211, y => 44),
  (x => 202, y => 45),
  (x => 203, y => 45),
  (x => 204, y => 45),
  (x => 205, y => 45),
  (x => 206, y => 45),
  (x => 207, y => 45),
  (x => 208, y => 45),
  (x => 209, y => 45),
  (x => 210, y => 45),
  (x => 204, y => 46),
  (x => 205, y => 46),
  (x => 206, y => 46),
  (x => 207, y => 46),
  (x => 208, y => 46),
  (x => 209, y => 46)
);
constant p1_9: CoordPairArray(0 to 182) := (
  (x => 203, y => 27),
  (x => 204, y => 27),
  (x => 205, y => 27),
  (x => 206, y => 27),
  (x => 207, y => 27),
  (x => 208, y => 27),
  (x => 201, y => 28),
  (x => 202, y => 28),
  (x => 203, y => 28),
  (x => 204, y => 28),
  (x => 205, y => 28),
  (x => 206, y => 28),
  (x => 207, y => 28),
  (x => 208, y => 28),
  (x => 209, y => 28),
  (x => 201, y => 29),
  (x => 202, y => 29),
  (x => 203, y => 29),
  (x => 204, y => 29),
  (x => 205, y => 29),
  (x => 206, y => 29),
  (x => 207, y => 29),
  (x => 208, y => 29),
  (x => 209, y => 29),
  (x => 200, y => 30),
  (x => 201, y => 30),
  (x => 202, y => 30),
  (x => 203, y => 30),
  (x => 204, y => 30),
  (x => 205, y => 30),
  (x => 206, y => 30),
  (x => 207, y => 30),
  (x => 208, y => 30),
  (x => 209, y => 30),
  (x => 210, y => 30),
  (x => 200, y => 31),
  (x => 201, y => 31),
  (x => 202, y => 31),
  (x => 203, y => 31),
  (x => 207, y => 31),
  (x => 208, y => 31),
  (x => 209, y => 31),
  (x => 210, y => 31),
  (x => 200, y => 32),
  (x => 201, y => 32),
  (x => 202, y => 32),
  (x => 203, y => 32),
  (x => 208, y => 32),
  (x => 209, y => 32),
  (x => 210, y => 32),
  (x => 211, y => 32),
  (x => 200, y => 33),
  (x => 201, y => 33),
  (x => 202, y => 33),
  (x => 208, y => 33),
  (x => 209, y => 33),
  (x => 210, y => 33),
  (x => 211, y => 33),
  (x => 199, y => 34),
  (x => 200, y => 34),
  (x => 201, y => 34),
  (x => 202, y => 34),
  (x => 208, y => 34),
  (x => 209, y => 34),
  (x => 210, y => 34),
  (x => 211, y => 34),
  (x => 199, y => 35),
  (x => 200, y => 35),
  (x => 201, y => 35),
  (x => 202, y => 35),
  (x => 208, y => 35),
  (x => 209, y => 35),
  (x => 210, y => 35),
  (x => 211, y => 35),
  (x => 200, y => 36),
  (x => 201, y => 36),
  (x => 202, y => 36),
  (x => 203, y => 36),
  (x => 208, y => 36),
  (x => 209, y => 36),
  (x => 210, y => 36),
  (x => 211, y => 36),
  (x => 200, y => 37),
  (x => 201, y => 37),
  (x => 202, y => 37),
  (x => 203, y => 37),
  (x => 207, y => 37),
  (x => 208, y => 37),
  (x => 209, y => 37),
  (x => 210, y => 37),
  (x => 211, y => 37),
  (x => 200, y => 38),
  (x => 201, y => 38),
  (x => 202, y => 38),
  (x => 203, y => 38),
  (x => 204, y => 38),
  (x => 205, y => 38),
  (x => 206, y => 38),
  (x => 207, y => 38),
  (x => 208, y => 38),
  (x => 209, y => 38),
  (x => 210, y => 38),
  (x => 211, y => 38),
  (x => 200, y => 39),
  (x => 201, y => 39),
  (x => 202, y => 39),
  (x => 203, y => 39),
  (x => 204, y => 39),
  (x => 205, y => 39),
  (x => 206, y => 39),
  (x => 207, y => 39),
  (x => 208, y => 39),
  (x => 209, y => 39),
  (x => 210, y => 39),
  (x => 211, y => 39),
  (x => 201, y => 40),
  (x => 202, y => 40),
  (x => 203, y => 40),
  (x => 204, y => 40),
  (x => 205, y => 40),
  (x => 208, y => 40),
  (x => 209, y => 40),
  (x => 210, y => 40),
  (x => 211, y => 40),
  (x => 203, y => 41),
  (x => 204, y => 41),
  (x => 208, y => 41),
  (x => 209, y => 41),
  (x => 210, y => 41),
  (x => 211, y => 41),
  (x => 208, y => 42),
  (x => 209, y => 42),
  (x => 210, y => 42),
  (x => 211, y => 42),
  (x => 208, y => 43),
  (x => 209, y => 43),
  (x => 210, y => 43),
  (x => 211, y => 43),
  (x => 207, y => 44),
  (x => 208, y => 44),
  (x => 209, y => 44),
  (x => 210, y => 44),
  (x => 207, y => 45),
  (x => 208, y => 45),
  (x => 209, y => 45),
  (x => 210, y => 45),
  (x => 206, y => 46),
  (x => 207, y => 46),
  (x => 208, y => 46),
  (x => 209, y => 46),
  (x => 210, y => 46),
  (x => 201, y => 47),
  (x => 202, y => 47),
  (x => 203, y => 47),
  (x => 204, y => 47),
  (x => 205, y => 47),
  (x => 206, y => 47),
  (x => 207, y => 47),
  (x => 208, y => 47),
  (x => 209, y => 47),
  (x => 201, y => 48),
  (x => 202, y => 48),
  (x => 203, y => 48),
  (x => 204, y => 48),
  (x => 205, y => 48),
  (x => 206, y => 48),
  (x => 207, y => 48),
  (x => 208, y => 48),
  (x => 209, y => 48),
  (x => 201, y => 49),
  (x => 202, y => 49),
  (x => 203, y => 49),
  (x => 204, y => 49),
  (x => 205, y => 49),
  (x => 206, y => 49),
  (x => 207, y => 49),
  (x => 208, y => 49),
  (x => 201, y => 50),
  (x => 202, y => 50),
  (x => 203, y => 50),
  (x => 204, y => 50),
  (x => 205, y => 50),
  (x => 206, y => 50)
);
constant p2_1: CoordPairArray(0 to 114) := (
  (x => 421, y => 26),
  (x => 422, y => 26),
  (x => 423, y => 26),
  (x => 420, y => 27),
  (x => 421, y => 27),
  (x => 422, y => 27),
  (x => 423, y => 27),
  (x => 418, y => 28),
  (x => 419, y => 28),
  (x => 420, y => 28),
  (x => 421, y => 28),
  (x => 422, y => 28),
  (x => 423, y => 28),
  (x => 416, y => 29),
  (x => 417, y => 29),
  (x => 418, y => 29),
  (x => 419, y => 29),
  (x => 420, y => 29),
  (x => 421, y => 29),
  (x => 422, y => 29),
  (x => 423, y => 29),
  (x => 415, y => 30),
  (x => 416, y => 30),
  (x => 417, y => 30),
  (x => 418, y => 30),
  (x => 419, y => 30),
  (x => 420, y => 30),
  (x => 421, y => 30),
  (x => 422, y => 30),
  (x => 423, y => 30),
  (x => 415, y => 31),
  (x => 416, y => 31),
  (x => 417, y => 31),
  (x => 418, y => 31),
  (x => 419, y => 31),
  (x => 420, y => 31),
  (x => 421, y => 31),
  (x => 422, y => 31),
  (x => 423, y => 31),
  (x => 415, y => 32),
  (x => 416, y => 32),
  (x => 417, y => 32),
  (x => 420, y => 32),
  (x => 421, y => 32),
  (x => 422, y => 32),
  (x => 423, y => 32),
  (x => 415, y => 33),
  (x => 420, y => 33),
  (x => 421, y => 33),
  (x => 422, y => 33),
  (x => 423, y => 33),
  (x => 420, y => 34),
  (x => 421, y => 34),
  (x => 422, y => 34),
  (x => 423, y => 34),
  (x => 420, y => 35),
  (x => 421, y => 35),
  (x => 422, y => 35),
  (x => 423, y => 35),
  (x => 420, y => 36),
  (x => 421, y => 36),
  (x => 422, y => 36),
  (x => 423, y => 36),
  (x => 420, y => 37),
  (x => 421, y => 37),
  (x => 422, y => 37),
  (x => 423, y => 37),
  (x => 420, y => 38),
  (x => 421, y => 38),
  (x => 422, y => 38),
  (x => 423, y => 38),
  (x => 420, y => 39),
  (x => 421, y => 39),
  (x => 422, y => 39),
  (x => 423, y => 39),
  (x => 420, y => 40),
  (x => 421, y => 40),
  (x => 422, y => 40),
  (x => 423, y => 40),
  (x => 420, y => 41),
  (x => 421, y => 41),
  (x => 422, y => 41),
  (x => 423, y => 41),
  (x => 420, y => 42),
  (x => 421, y => 42),
  (x => 422, y => 42),
  (x => 423, y => 42),
  (x => 420, y => 43),
  (x => 421, y => 43),
  (x => 422, y => 43),
  (x => 423, y => 43),
  (x => 420, y => 44),
  (x => 421, y => 44),
  (x => 422, y => 44),
  (x => 423, y => 44),
  (x => 420, y => 45),
  (x => 421, y => 45),
  (x => 422, y => 45),
  (x => 423, y => 45),
  (x => 420, y => 46),
  (x => 421, y => 46),
  (x => 422, y => 46),
  (x => 423, y => 46),
  (x => 420, y => 47),
  (x => 421, y => 47),
  (x => 422, y => 47),
  (x => 423, y => 47),
  (x => 420, y => 48),
  (x => 421, y => 48),
  (x => 422, y => 48),
  (x => 423, y => 48),
  (x => 420, y => 49),
  (x => 421, y => 49),
  (x => 422, y => 49),
  (x => 423, y => 49)
);
constant p2_2: CoordPairArray(0 to 157) := (
  (x => 419, y => 23),
  (x => 420, y => 23),
  (x => 421, y => 23),
  (x => 422, y => 23),
  (x => 416, y => 24),
  (x => 417, y => 24),
  (x => 418, y => 24),
  (x => 419, y => 24),
  (x => 420, y => 24),
  (x => 421, y => 24),
  (x => 422, y => 24),
  (x => 423, y => 24),
  (x => 424, y => 24),
  (x => 416, y => 25),
  (x => 417, y => 25),
  (x => 418, y => 25),
  (x => 419, y => 25),
  (x => 420, y => 25),
  (x => 421, y => 25),
  (x => 422, y => 25),
  (x => 423, y => 25),
  (x => 424, y => 25),
  (x => 425, y => 25),
  (x => 416, y => 26),
  (x => 417, y => 26),
  (x => 418, y => 26),
  (x => 419, y => 26),
  (x => 420, y => 26),
  (x => 421, y => 26),
  (x => 422, y => 26),
  (x => 423, y => 26),
  (x => 424, y => 26),
  (x => 425, y => 26),
  (x => 416, y => 27),
  (x => 417, y => 27),
  (x => 418, y => 27),
  (x => 419, y => 27),
  (x => 420, y => 27),
  (x => 421, y => 27),
  (x => 422, y => 27),
  (x => 423, y => 27),
  (x => 424, y => 27),
  (x => 425, y => 27),
  (x => 426, y => 27),
  (x => 416, y => 28),
  (x => 422, y => 28),
  (x => 423, y => 28),
  (x => 424, y => 28),
  (x => 425, y => 28),
  (x => 426, y => 28),
  (x => 423, y => 29),
  (x => 424, y => 29),
  (x => 425, y => 29),
  (x => 426, y => 29),
  (x => 423, y => 30),
  (x => 424, y => 30),
  (x => 425, y => 30),
  (x => 426, y => 30),
  (x => 423, y => 31),
  (x => 424, y => 31),
  (x => 425, y => 31),
  (x => 426, y => 31),
  (x => 423, y => 32),
  (x => 424, y => 32),
  (x => 425, y => 32),
  (x => 426, y => 32),
  (x => 422, y => 33),
  (x => 423, y => 33),
  (x => 424, y => 33),
  (x => 425, y => 33),
  (x => 421, y => 34),
  (x => 422, y => 34),
  (x => 423, y => 34),
  (x => 424, y => 34),
  (x => 425, y => 34),
  (x => 420, y => 35),
  (x => 421, y => 35),
  (x => 422, y => 35),
  (x => 423, y => 35),
  (x => 424, y => 35),
  (x => 419, y => 36),
  (x => 420, y => 36),
  (x => 421, y => 36),
  (x => 422, y => 36),
  (x => 423, y => 36),
  (x => 418, y => 37),
  (x => 419, y => 37),
  (x => 420, y => 37),
  (x => 421, y => 37),
  (x => 422, y => 37),
  (x => 418, y => 38),
  (x => 419, y => 38),
  (x => 420, y => 38),
  (x => 421, y => 38),
  (x => 417, y => 39),
  (x => 418, y => 39),
  (x => 419, y => 39),
  (x => 420, y => 39),
  (x => 416, y => 40),
  (x => 417, y => 40),
  (x => 418, y => 40),
  (x => 419, y => 40),
  (x => 416, y => 41),
  (x => 417, y => 41),
  (x => 418, y => 41),
  (x => 419, y => 41),
  (x => 416, y => 42),
  (x => 417, y => 42),
  (x => 418, y => 42),
  (x => 419, y => 42),
  (x => 415, y => 43),
  (x => 416, y => 43),
  (x => 417, y => 43),
  (x => 418, y => 43),
  (x => 419, y => 43),
  (x => 420, y => 43),
  (x => 421, y => 43),
  (x => 422, y => 43),
  (x => 423, y => 43),
  (x => 424, y => 43),
  (x => 425, y => 43),
  (x => 426, y => 43),
  (x => 415, y => 44),
  (x => 416, y => 44),
  (x => 417, y => 44),
  (x => 418, y => 44),
  (x => 419, y => 44),
  (x => 420, y => 44),
  (x => 421, y => 44),
  (x => 422, y => 44),
  (x => 423, y => 44),
  (x => 424, y => 44),
  (x => 425, y => 44),
  (x => 426, y => 44),
  (x => 415, y => 45),
  (x => 416, y => 45),
  (x => 417, y => 45),
  (x => 418, y => 45),
  (x => 419, y => 45),
  (x => 420, y => 45),
  (x => 421, y => 45),
  (x => 422, y => 45),
  (x => 423, y => 45),
  (x => 424, y => 45),
  (x => 425, y => 45),
  (x => 426, y => 45),
  (x => 415, y => 46),
  (x => 416, y => 46),
  (x => 417, y => 46),
  (x => 418, y => 46),
  (x => 419, y => 46),
  (x => 420, y => 46),
  (x => 421, y => 46),
  (x => 422, y => 46),
  (x => 423, y => 46),
  (x => 424, y => 46),
  (x => 425, y => 46),
  (x => 426, y => 46)
);
constant p2_3: CoordPairArray(0 to 151) := (
  (x => 418, y => 22),
  (x => 419, y => 22),
  (x => 420, y => 22),
  (x => 421, y => 22),
  (x => 422, y => 22),
  (x => 416, y => 23),
  (x => 417, y => 23),
  (x => 418, y => 23),
  (x => 419, y => 23),
  (x => 420, y => 23),
  (x => 421, y => 23),
  (x => 422, y => 23),
  (x => 423, y => 23),
  (x => 424, y => 23),
  (x => 416, y => 24),
  (x => 417, y => 24),
  (x => 418, y => 24),
  (x => 419, y => 24),
  (x => 420, y => 24),
  (x => 421, y => 24),
  (x => 422, y => 24),
  (x => 423, y => 24),
  (x => 424, y => 24),
  (x => 425, y => 24),
  (x => 416, y => 25),
  (x => 417, y => 25),
  (x => 418, y => 25),
  (x => 419, y => 25),
  (x => 420, y => 25),
  (x => 421, y => 25),
  (x => 422, y => 25),
  (x => 423, y => 25),
  (x => 424, y => 25),
  (x => 425, y => 25),
  (x => 416, y => 26),
  (x => 421, y => 26),
  (x => 422, y => 26),
  (x => 423, y => 26),
  (x => 424, y => 26),
  (x => 425, y => 26),
  (x => 422, y => 27),
  (x => 423, y => 27),
  (x => 424, y => 27),
  (x => 425, y => 27),
  (x => 422, y => 28),
  (x => 423, y => 28),
  (x => 424, y => 28),
  (x => 425, y => 28),
  (x => 422, y => 29),
  (x => 423, y => 29),
  (x => 424, y => 29),
  (x => 425, y => 29),
  (x => 422, y => 30),
  (x => 423, y => 30),
  (x => 424, y => 30),
  (x => 425, y => 30),
  (x => 421, y => 31),
  (x => 422, y => 31),
  (x => 423, y => 31),
  (x => 424, y => 31),
  (x => 417, y => 32),
  (x => 418, y => 32),
  (x => 419, y => 32),
  (x => 420, y => 32),
  (x => 421, y => 32),
  (x => 422, y => 32),
  (x => 423, y => 32),
  (x => 424, y => 32),
  (x => 418, y => 33),
  (x => 419, y => 33),
  (x => 420, y => 33),
  (x => 421, y => 33),
  (x => 422, y => 33),
  (x => 418, y => 34),
  (x => 419, y => 34),
  (x => 420, y => 34),
  (x => 421, y => 34),
  (x => 422, y => 34),
  (x => 417, y => 35),
  (x => 418, y => 35),
  (x => 419, y => 35),
  (x => 420, y => 35),
  (x => 421, y => 35),
  (x => 422, y => 35),
  (x => 423, y => 35),
  (x => 424, y => 35),
  (x => 421, y => 36),
  (x => 422, y => 36),
  (x => 423, y => 36),
  (x => 424, y => 36),
  (x => 425, y => 36),
  (x => 422, y => 37),
  (x => 423, y => 37),
  (x => 424, y => 37),
  (x => 425, y => 37),
  (x => 423, y => 38),
  (x => 424, y => 38),
  (x => 425, y => 38),
  (x => 426, y => 38),
  (x => 423, y => 39),
  (x => 424, y => 39),
  (x => 425, y => 39),
  (x => 426, y => 39),
  (x => 423, y => 40),
  (x => 424, y => 40),
  (x => 425, y => 40),
  (x => 426, y => 40),
  (x => 422, y => 41),
  (x => 423, y => 41),
  (x => 424, y => 41),
  (x => 425, y => 41),
  (x => 426, y => 41),
  (x => 416, y => 42),
  (x => 417, y => 42),
  (x => 420, y => 42),
  (x => 421, y => 42),
  (x => 422, y => 42),
  (x => 423, y => 42),
  (x => 424, y => 42),
  (x => 425, y => 42),
  (x => 416, y => 43),
  (x => 417, y => 43),
  (x => 418, y => 43),
  (x => 419, y => 43),
  (x => 420, y => 43),
  (x => 421, y => 43),
  (x => 422, y => 43),
  (x => 423, y => 43),
  (x => 424, y => 43),
  (x => 425, y => 43),
  (x => 416, y => 44),
  (x => 417, y => 44),
  (x => 418, y => 44),
  (x => 419, y => 44),
  (x => 420, y => 44),
  (x => 421, y => 44),
  (x => 422, y => 44),
  (x => 423, y => 44),
  (x => 424, y => 44),
  (x => 415, y => 45),
  (x => 416, y => 45),
  (x => 417, y => 45),
  (x => 418, y => 45),
  (x => 419, y => 45),
  (x => 420, y => 45),
  (x => 421, y => 45),
  (x => 422, y => 45),
  (x => 423, y => 45),
  (x => 418, y => 46),
  (x => 419, y => 46),
  (x => 420, y => 46),
  (x => 421, y => 46)
);
constant p2_4: CoordPairArray(0 to 173) := (
  (x => 419, y => 20),
  (x => 420, y => 20),
  (x => 421, y => 20),
  (x => 422, y => 20),
  (x => 423, y => 20),
  (x => 419, y => 21),
  (x => 420, y => 21),
  (x => 421, y => 21),
  (x => 422, y => 21),
  (x => 423, y => 21),
  (x => 419, y => 22),
  (x => 420, y => 22),
  (x => 421, y => 22),
  (x => 422, y => 22),
  (x => 423, y => 22),
  (x => 418, y => 23),
  (x => 419, y => 23),
  (x => 420, y => 23),
  (x => 421, y => 23),
  (x => 422, y => 23),
  (x => 423, y => 23),
  (x => 418, y => 24),
  (x => 419, y => 24),
  (x => 420, y => 24),
  (x => 421, y => 24),
  (x => 422, y => 24),
  (x => 423, y => 24),
  (x => 417, y => 25),
  (x => 418, y => 25),
  (x => 419, y => 25),
  (x => 420, y => 25),
  (x => 421, y => 25),
  (x => 422, y => 25),
  (x => 423, y => 25),
  (x => 417, y => 26),
  (x => 418, y => 26),
  (x => 419, y => 26),
  (x => 420, y => 26),
  (x => 421, y => 26),
  (x => 422, y => 26),
  (x => 423, y => 26),
  (x => 416, y => 27),
  (x => 417, y => 27),
  (x => 418, y => 27),
  (x => 420, y => 27),
  (x => 421, y => 27),
  (x => 422, y => 27),
  (x => 423, y => 27),
  (x => 416, y => 28),
  (x => 417, y => 28),
  (x => 420, y => 28),
  (x => 421, y => 28),
  (x => 422, y => 28),
  (x => 423, y => 28),
  (x => 415, y => 29),
  (x => 416, y => 29),
  (x => 417, y => 29),
  (x => 420, y => 29),
  (x => 421, y => 29),
  (x => 422, y => 29),
  (x => 423, y => 29),
  (x => 415, y => 30),
  (x => 416, y => 30),
  (x => 417, y => 30),
  (x => 420, y => 30),
  (x => 421, y => 30),
  (x => 422, y => 30),
  (x => 423, y => 30),
  (x => 414, y => 31),
  (x => 415, y => 31),
  (x => 416, y => 31),
  (x => 420, y => 31),
  (x => 421, y => 31),
  (x => 422, y => 31),
  (x => 423, y => 31),
  (x => 414, y => 32),
  (x => 415, y => 32),
  (x => 416, y => 32),
  (x => 420, y => 32),
  (x => 421, y => 32),
  (x => 422, y => 32),
  (x => 423, y => 32),
  (x => 413, y => 33),
  (x => 414, y => 33),
  (x => 415, y => 33),
  (x => 420, y => 33),
  (x => 421, y => 33),
  (x => 422, y => 33),
  (x => 423, y => 33),
  (x => 413, y => 34),
  (x => 414, y => 34),
  (x => 420, y => 34),
  (x => 421, y => 34),
  (x => 422, y => 34),
  (x => 423, y => 34),
  (x => 412, y => 35),
  (x => 413, y => 35),
  (x => 414, y => 35),
  (x => 420, y => 35),
  (x => 421, y => 35),
  (x => 422, y => 35),
  (x => 423, y => 35),
  (x => 412, y => 36),
  (x => 413, y => 36),
  (x => 414, y => 36),
  (x => 415, y => 36),
  (x => 416, y => 36),
  (x => 417, y => 36),
  (x => 418, y => 36),
  (x => 419, y => 36),
  (x => 420, y => 36),
  (x => 421, y => 36),
  (x => 422, y => 36),
  (x => 423, y => 36),
  (x => 424, y => 36),
  (x => 425, y => 36),
  (x => 412, y => 37),
  (x => 413, y => 37),
  (x => 414, y => 37),
  (x => 415, y => 37),
  (x => 416, y => 37),
  (x => 417, y => 37),
  (x => 418, y => 37),
  (x => 419, y => 37),
  (x => 420, y => 37),
  (x => 421, y => 37),
  (x => 422, y => 37),
  (x => 423, y => 37),
  (x => 424, y => 37),
  (x => 425, y => 37),
  (x => 412, y => 38),
  (x => 413, y => 38),
  (x => 414, y => 38),
  (x => 415, y => 38),
  (x => 416, y => 38),
  (x => 417, y => 38),
  (x => 418, y => 38),
  (x => 419, y => 38),
  (x => 420, y => 38),
  (x => 421, y => 38),
  (x => 422, y => 38),
  (x => 423, y => 38),
  (x => 424, y => 38),
  (x => 425, y => 38),
  (x => 412, y => 39),
  (x => 413, y => 39),
  (x => 414, y => 39),
  (x => 415, y => 39),
  (x => 416, y => 39),
  (x => 417, y => 39),
  (x => 418, y => 39),
  (x => 419, y => 39),
  (x => 420, y => 39),
  (x => 421, y => 39),
  (x => 422, y => 39),
  (x => 423, y => 39),
  (x => 424, y => 39),
  (x => 425, y => 39),
  (x => 420, y => 40),
  (x => 421, y => 40),
  (x => 422, y => 40),
  (x => 423, y => 40),
  (x => 420, y => 41),
  (x => 421, y => 41),
  (x => 422, y => 41),
  (x => 423, y => 41),
  (x => 420, y => 42),
  (x => 421, y => 42),
  (x => 422, y => 42),
  (x => 423, y => 42),
  (x => 420, y => 43),
  (x => 421, y => 43),
  (x => 422, y => 43),
  (x => 423, y => 43)
);
constant p2_5: CoordPairArray(0 to 158) := (
  (x => 420, y => 23),
  (x => 421, y => 23),
  (x => 422, y => 23),
  (x => 423, y => 23),
  (x => 424, y => 23),
  (x => 425, y => 23),
  (x => 426, y => 23),
  (x => 427, y => 23),
  (x => 428, y => 23),
  (x => 420, y => 24),
  (x => 421, y => 24),
  (x => 422, y => 24),
  (x => 423, y => 24),
  (x => 424, y => 24),
  (x => 425, y => 24),
  (x => 426, y => 24),
  (x => 427, y => 24),
  (x => 428, y => 24),
  (x => 420, y => 25),
  (x => 421, y => 25),
  (x => 422, y => 25),
  (x => 423, y => 25),
  (x => 424, y => 25),
  (x => 425, y => 25),
  (x => 426, y => 25),
  (x => 427, y => 25),
  (x => 428, y => 25),
  (x => 420, y => 26),
  (x => 421, y => 26),
  (x => 422, y => 26),
  (x => 423, y => 26),
  (x => 424, y => 26),
  (x => 425, y => 26),
  (x => 426, y => 26),
  (x => 427, y => 26),
  (x => 428, y => 26),
  (x => 420, y => 27),
  (x => 421, y => 27),
  (x => 422, y => 27),
  (x => 420, y => 28),
  (x => 421, y => 28),
  (x => 422, y => 28),
  (x => 420, y => 29),
  (x => 421, y => 29),
  (x => 422, y => 29),
  (x => 419, y => 30),
  (x => 420, y => 30),
  (x => 421, y => 30),
  (x => 422, y => 30),
  (x => 419, y => 31),
  (x => 420, y => 31),
  (x => 421, y => 31),
  (x => 419, y => 32),
  (x => 420, y => 32),
  (x => 421, y => 32),
  (x => 422, y => 32),
  (x => 423, y => 32),
  (x => 424, y => 32),
  (x => 425, y => 32),
  (x => 426, y => 32),
  (x => 427, y => 32),
  (x => 419, y => 33),
  (x => 420, y => 33),
  (x => 421, y => 33),
  (x => 422, y => 33),
  (x => 423, y => 33),
  (x => 424, y => 33),
  (x => 425, y => 33),
  (x => 426, y => 33),
  (x => 427, y => 33),
  (x => 428, y => 33),
  (x => 419, y => 34),
  (x => 420, y => 34),
  (x => 421, y => 34),
  (x => 422, y => 34),
  (x => 423, y => 34),
  (x => 424, y => 34),
  (x => 425, y => 34),
  (x => 426, y => 34),
  (x => 427, y => 34),
  (x => 428, y => 34),
  (x => 419, y => 35),
  (x => 420, y => 35),
  (x => 421, y => 35),
  (x => 422, y => 35),
  (x => 423, y => 35),
  (x => 424, y => 35),
  (x => 425, y => 35),
  (x => 426, y => 35),
  (x => 427, y => 35),
  (x => 428, y => 35),
  (x => 429, y => 35),
  (x => 424, y => 36),
  (x => 425, y => 36),
  (x => 426, y => 36),
  (x => 427, y => 36),
  (x => 428, y => 36),
  (x => 429, y => 36),
  (x => 425, y => 37),
  (x => 426, y => 37),
  (x => 427, y => 37),
  (x => 428, y => 37),
  (x => 429, y => 37),
  (x => 426, y => 38),
  (x => 427, y => 38),
  (x => 428, y => 38),
  (x => 429, y => 38),
  (x => 426, y => 39),
  (x => 427, y => 39),
  (x => 428, y => 39),
  (x => 429, y => 39),
  (x => 426, y => 40),
  (x => 427, y => 40),
  (x => 428, y => 40),
  (x => 429, y => 40),
  (x => 425, y => 41),
  (x => 426, y => 41),
  (x => 427, y => 41),
  (x => 428, y => 41),
  (x => 429, y => 41),
  (x => 419, y => 42),
  (x => 420, y => 42),
  (x => 423, y => 42),
  (x => 424, y => 42),
  (x => 425, y => 42),
  (x => 426, y => 42),
  (x => 427, y => 42),
  (x => 428, y => 42),
  (x => 419, y => 43),
  (x => 420, y => 43),
  (x => 421, y => 43),
  (x => 422, y => 43),
  (x => 423, y => 43),
  (x => 424, y => 43),
  (x => 425, y => 43),
  (x => 426, y => 43),
  (x => 427, y => 43),
  (x => 428, y => 43),
  (x => 419, y => 44),
  (x => 420, y => 44),
  (x => 421, y => 44),
  (x => 422, y => 44),
  (x => 423, y => 44),
  (x => 424, y => 44),
  (x => 425, y => 44),
  (x => 426, y => 44),
  (x => 427, y => 44),
  (x => 419, y => 45),
  (x => 420, y => 45),
  (x => 421, y => 45),
  (x => 422, y => 45),
  (x => 423, y => 45),
  (x => 424, y => 45),
  (x => 425, y => 45),
  (x => 426, y => 45),
  (x => 421, y => 46),
  (x => 422, y => 46),
  (x => 423, y => 46),
  (x => 424, y => 46)
);
constant p2_6: CoordPairArray(0 to 185) := (
  (x => 426, y => 20),
  (x => 427, y => 20),
  (x => 428, y => 20),
  (x => 429, y => 20),
  (x => 430, y => 20),
  (x => 431, y => 20),
  (x => 424, y => 21),
  (x => 425, y => 21),
  (x => 426, y => 21),
  (x => 427, y => 21),
  (x => 428, y => 21),
  (x => 429, y => 21),
  (x => 430, y => 21),
  (x => 431, y => 21),
  (x => 423, y => 22),
  (x => 424, y => 22),
  (x => 425, y => 22),
  (x => 426, y => 22),
  (x => 427, y => 22),
  (x => 428, y => 22),
  (x => 429, y => 22),
  (x => 430, y => 22),
  (x => 431, y => 22),
  (x => 423, y => 23),
  (x => 424, y => 23),
  (x => 425, y => 23),
  (x => 426, y => 23),
  (x => 427, y => 23),
  (x => 428, y => 23),
  (x => 429, y => 23),
  (x => 430, y => 23),
  (x => 431, y => 23),
  (x => 422, y => 24),
  (x => 423, y => 24),
  (x => 424, y => 24),
  (x => 425, y => 24),
  (x => 426, y => 24),
  (x => 422, y => 25),
  (x => 423, y => 25),
  (x => 424, y => 25),
  (x => 425, y => 25),
  (x => 421, y => 26),
  (x => 422, y => 26),
  (x => 423, y => 26),
  (x => 424, y => 26),
  (x => 421, y => 27),
  (x => 422, y => 27),
  (x => 423, y => 27),
  (x => 424, y => 27),
  (x => 421, y => 28),
  (x => 422, y => 28),
  (x => 423, y => 28),
  (x => 424, y => 28),
  (x => 421, y => 29),
  (x => 422, y => 29),
  (x => 423, y => 29),
  (x => 427, y => 29),
  (x => 428, y => 29),
  (x => 429, y => 29),
  (x => 430, y => 29),
  (x => 421, y => 30),
  (x => 422, y => 30),
  (x => 423, y => 30),
  (x => 424, y => 30),
  (x => 425, y => 30),
  (x => 426, y => 30),
  (x => 427, y => 30),
  (x => 428, y => 30),
  (x => 429, y => 30),
  (x => 430, y => 30),
  (x => 431, y => 30),
  (x => 421, y => 31),
  (x => 422, y => 31),
  (x => 423, y => 31),
  (x => 424, y => 31),
  (x => 425, y => 31),
  (x => 426, y => 31),
  (x => 427, y => 31),
  (x => 428, y => 31),
  (x => 429, y => 31),
  (x => 430, y => 31),
  (x => 431, y => 31),
  (x => 421, y => 32),
  (x => 422, y => 32),
  (x => 423, y => 32),
  (x => 424, y => 32),
  (x => 425, y => 32),
  (x => 426, y => 32),
  (x => 427, y => 32),
  (x => 428, y => 32),
  (x => 429, y => 32),
  (x => 430, y => 32),
  (x => 431, y => 32),
  (x => 432, y => 32),
  (x => 421, y => 33),
  (x => 422, y => 33),
  (x => 423, y => 33),
  (x => 424, y => 33),
  (x => 429, y => 33),
  (x => 430, y => 33),
  (x => 431, y => 33),
  (x => 432, y => 33),
  (x => 421, y => 34),
  (x => 422, y => 34),
  (x => 423, y => 34),
  (x => 424, y => 34),
  (x => 429, y => 34),
  (x => 430, y => 34),
  (x => 431, y => 34),
  (x => 432, y => 34),
  (x => 421, y => 35),
  (x => 422, y => 35),
  (x => 423, y => 35),
  (x => 424, y => 35),
  (x => 429, y => 35),
  (x => 430, y => 35),
  (x => 431, y => 35),
  (x => 432, y => 35),
  (x => 421, y => 36),
  (x => 422, y => 36),
  (x => 423, y => 36),
  (x => 424, y => 36),
  (x => 429, y => 36),
  (x => 430, y => 36),
  (x => 431, y => 36),
  (x => 432, y => 36),
  (x => 421, y => 37),
  (x => 422, y => 37),
  (x => 423, y => 37),
  (x => 424, y => 37),
  (x => 429, y => 37),
  (x => 430, y => 37),
  (x => 431, y => 37),
  (x => 432, y => 37),
  (x => 421, y => 38),
  (x => 422, y => 38),
  (x => 423, y => 38),
  (x => 424, y => 38),
  (x => 429, y => 38),
  (x => 430, y => 38),
  (x => 431, y => 38),
  (x => 432, y => 38),
  (x => 421, y => 39),
  (x => 422, y => 39),
  (x => 423, y => 39),
  (x => 424, y => 39),
  (x => 425, y => 39),
  (x => 428, y => 39),
  (x => 429, y => 39),
  (x => 430, y => 39),
  (x => 431, y => 39),
  (x => 432, y => 39),
  (x => 422, y => 40),
  (x => 423, y => 40),
  (x => 424, y => 40),
  (x => 425, y => 40),
  (x => 426, y => 40),
  (x => 427, y => 40),
  (x => 428, y => 40),
  (x => 429, y => 40),
  (x => 430, y => 40),
  (x => 431, y => 40),
  (x => 422, y => 41),
  (x => 423, y => 41),
  (x => 424, y => 41),
  (x => 425, y => 41),
  (x => 426, y => 41),
  (x => 427, y => 41),
  (x => 428, y => 41),
  (x => 429, y => 41),
  (x => 430, y => 41),
  (x => 431, y => 41),
  (x => 423, y => 42),
  (x => 424, y => 42),
  (x => 425, y => 42),
  (x => 426, y => 42),
  (x => 427, y => 42),
  (x => 428, y => 42),
  (x => 429, y => 42),
  (x => 430, y => 42),
  (x => 424, y => 43),
  (x => 425, y => 43),
  (x => 426, y => 43),
  (x => 427, y => 43),
  (x => 428, y => 43),
  (x => 429, y => 43)
);
constant p2_7: CoordPairArray(0 to 135) := (
  (x => 426, y => 23),
  (x => 427, y => 23),
  (x => 428, y => 23),
  (x => 429, y => 23),
  (x => 430, y => 23),
  (x => 431, y => 23),
  (x => 432, y => 23),
  (x => 433, y => 23),
  (x => 434, y => 23),
  (x => 435, y => 23),
  (x => 436, y => 23),
  (x => 437, y => 23),
  (x => 426, y => 24),
  (x => 427, y => 24),
  (x => 428, y => 24),
  (x => 429, y => 24),
  (x => 430, y => 24),
  (x => 431, y => 24),
  (x => 432, y => 24),
  (x => 433, y => 24),
  (x => 434, y => 24),
  (x => 435, y => 24),
  (x => 436, y => 24),
  (x => 437, y => 24),
  (x => 426, y => 25),
  (x => 427, y => 25),
  (x => 428, y => 25),
  (x => 429, y => 25),
  (x => 430, y => 25),
  (x => 431, y => 25),
  (x => 432, y => 25),
  (x => 433, y => 25),
  (x => 434, y => 25),
  (x => 435, y => 25),
  (x => 436, y => 25),
  (x => 437, y => 25),
  (x => 426, y => 26),
  (x => 427, y => 26),
  (x => 428, y => 26),
  (x => 429, y => 26),
  (x => 430, y => 26),
  (x => 431, y => 26),
  (x => 432, y => 26),
  (x => 433, y => 26),
  (x => 434, y => 26),
  (x => 435, y => 26),
  (x => 436, y => 26),
  (x => 437, y => 26),
  (x => 426, y => 27),
  (x => 427, y => 27),
  (x => 428, y => 27),
  (x => 429, y => 27),
  (x => 430, y => 27),
  (x => 431, y => 27),
  (x => 432, y => 27),
  (x => 433, y => 27),
  (x => 434, y => 27),
  (x => 435, y => 27),
  (x => 436, y => 27),
  (x => 437, y => 27),
  (x => 434, y => 28),
  (x => 435, y => 28),
  (x => 436, y => 28),
  (x => 434, y => 29),
  (x => 435, y => 29),
  (x => 436, y => 29),
  (x => 433, y => 30),
  (x => 434, y => 30),
  (x => 435, y => 30),
  (x => 436, y => 30),
  (x => 433, y => 31),
  (x => 434, y => 31),
  (x => 435, y => 31),
  (x => 432, y => 32),
  (x => 433, y => 32),
  (x => 434, y => 32),
  (x => 435, y => 32),
  (x => 432, y => 33),
  (x => 433, y => 33),
  (x => 434, y => 33),
  (x => 435, y => 33),
  (x => 431, y => 34),
  (x => 432, y => 34),
  (x => 433, y => 34),
  (x => 434, y => 34),
  (x => 431, y => 35),
  (x => 432, y => 35),
  (x => 433, y => 35),
  (x => 434, y => 35),
  (x => 431, y => 36),
  (x => 432, y => 36),
  (x => 433, y => 36),
  (x => 434, y => 36),
  (x => 430, y => 37),
  (x => 431, y => 37),
  (x => 432, y => 37),
  (x => 433, y => 37),
  (x => 430, y => 38),
  (x => 431, y => 38),
  (x => 432, y => 38),
  (x => 433, y => 38),
  (x => 430, y => 39),
  (x => 431, y => 39),
  (x => 432, y => 39),
  (x => 433, y => 39),
  (x => 429, y => 40),
  (x => 430, y => 40),
  (x => 431, y => 40),
  (x => 432, y => 40),
  (x => 433, y => 40),
  (x => 429, y => 41),
  (x => 430, y => 41),
  (x => 431, y => 41),
  (x => 432, y => 41),
  (x => 429, y => 42),
  (x => 430, y => 42),
  (x => 431, y => 42),
  (x => 432, y => 42),
  (x => 429, y => 43),
  (x => 430, y => 43),
  (x => 431, y => 43),
  (x => 432, y => 43),
  (x => 429, y => 44),
  (x => 430, y => 44),
  (x => 431, y => 44),
  (x => 432, y => 44),
  (x => 428, y => 45),
  (x => 429, y => 45),
  (x => 430, y => 45),
  (x => 431, y => 45),
  (x => 432, y => 45),
  (x => 428, y => 46),
  (x => 429, y => 46),
  (x => 430, y => 46),
  (x => 431, y => 46),
  (x => 432, y => 46)
);
constant p2_8: CoordPairArray(0 to 191) := (
  (x => 434, y => 20),
  (x => 435, y => 20),
  (x => 436, y => 20),
  (x => 437, y => 20),
  (x => 432, y => 21),
  (x => 433, y => 21),
  (x => 434, y => 21),
  (x => 435, y => 21),
  (x => 436, y => 21),
  (x => 437, y => 21),
  (x => 438, y => 21),
  (x => 439, y => 21),
  (x => 431, y => 22),
  (x => 432, y => 22),
  (x => 433, y => 22),
  (x => 434, y => 22),
  (x => 435, y => 22),
  (x => 436, y => 22),
  (x => 437, y => 22),
  (x => 438, y => 22),
  (x => 439, y => 22),
  (x => 440, y => 22),
  (x => 431, y => 23),
  (x => 432, y => 23),
  (x => 433, y => 23),
  (x => 434, y => 23),
  (x => 435, y => 23),
  (x => 436, y => 23),
  (x => 437, y => 23),
  (x => 438, y => 23),
  (x => 439, y => 23),
  (x => 440, y => 23),
  (x => 441, y => 23),
  (x => 430, y => 24),
  (x => 431, y => 24),
  (x => 432, y => 24),
  (x => 433, y => 24),
  (x => 438, y => 24),
  (x => 439, y => 24),
  (x => 440, y => 24),
  (x => 441, y => 24),
  (x => 430, y => 25),
  (x => 431, y => 25),
  (x => 432, y => 25),
  (x => 433, y => 25),
  (x => 438, y => 25),
  (x => 439, y => 25),
  (x => 440, y => 25),
  (x => 441, y => 25),
  (x => 430, y => 26),
  (x => 431, y => 26),
  (x => 432, y => 26),
  (x => 433, y => 26),
  (x => 439, y => 26),
  (x => 440, y => 26),
  (x => 441, y => 26),
  (x => 430, y => 27),
  (x => 431, y => 27),
  (x => 432, y => 27),
  (x => 433, y => 27),
  (x => 439, y => 27),
  (x => 440, y => 27),
  (x => 441, y => 27),
  (x => 430, y => 28),
  (x => 431, y => 28),
  (x => 432, y => 28),
  (x => 433, y => 28),
  (x => 438, y => 28),
  (x => 439, y => 28),
  (x => 440, y => 28),
  (x => 441, y => 28),
  (x => 431, y => 29),
  (x => 432, y => 29),
  (x => 433, y => 29),
  (x => 434, y => 29),
  (x => 438, y => 29),
  (x => 439, y => 29),
  (x => 440, y => 29),
  (x => 432, y => 30),
  (x => 433, y => 30),
  (x => 434, y => 30),
  (x => 435, y => 30),
  (x => 436, y => 30),
  (x => 437, y => 30),
  (x => 438, y => 30),
  (x => 439, y => 30),
  (x => 433, y => 31),
  (x => 434, y => 31),
  (x => 435, y => 31),
  (x => 436, y => 31),
  (x => 437, y => 31),
  (x => 438, y => 31),
  (x => 433, y => 32),
  (x => 434, y => 32),
  (x => 435, y => 32),
  (x => 436, y => 32),
  (x => 437, y => 32),
  (x => 438, y => 32),
  (x => 431, y => 33),
  (x => 432, y => 33),
  (x => 433, y => 33),
  (x => 434, y => 33),
  (x => 435, y => 33),
  (x => 436, y => 33),
  (x => 437, y => 33),
  (x => 438, y => 33),
  (x => 439, y => 33),
  (x => 440, y => 33),
  (x => 430, y => 34),
  (x => 431, y => 34),
  (x => 432, y => 34),
  (x => 433, y => 34),
  (x => 434, y => 34),
  (x => 437, y => 34),
  (x => 438, y => 34),
  (x => 439, y => 34),
  (x => 440, y => 34),
  (x => 441, y => 34),
  (x => 430, y => 35),
  (x => 431, y => 35),
  (x => 432, y => 35),
  (x => 433, y => 35),
  (x => 438, y => 35),
  (x => 439, y => 35),
  (x => 440, y => 35),
  (x => 441, y => 35),
  (x => 430, y => 36),
  (x => 431, y => 36),
  (x => 432, y => 36),
  (x => 439, y => 36),
  (x => 440, y => 36),
  (x => 441, y => 36),
  (x => 430, y => 37),
  (x => 431, y => 37),
  (x => 432, y => 37),
  (x => 439, y => 37),
  (x => 440, y => 37),
  (x => 441, y => 37),
  (x => 430, y => 38),
  (x => 431, y => 38),
  (x => 432, y => 38),
  (x => 439, y => 38),
  (x => 440, y => 38),
  (x => 441, y => 38),
  (x => 430, y => 39),
  (x => 431, y => 39),
  (x => 432, y => 39),
  (x => 439, y => 39),
  (x => 440, y => 39),
  (x => 441, y => 39),
  (x => 430, y => 40),
  (x => 431, y => 40),
  (x => 432, y => 40),
  (x => 433, y => 40),
  (x => 438, y => 40),
  (x => 439, y => 40),
  (x => 440, y => 40),
  (x => 441, y => 40),
  (x => 430, y => 41),
  (x => 431, y => 41),
  (x => 432, y => 41),
  (x => 433, y => 41),
  (x => 434, y => 41),
  (x => 435, y => 41),
  (x => 436, y => 41),
  (x => 437, y => 41),
  (x => 438, y => 41),
  (x => 439, y => 41),
  (x => 440, y => 41),
  (x => 441, y => 41),
  (x => 431, y => 42),
  (x => 432, y => 42),
  (x => 433, y => 42),
  (x => 434, y => 42),
  (x => 435, y => 42),
  (x => 436, y => 42),
  (x => 437, y => 42),
  (x => 438, y => 42),
  (x => 439, y => 42),
  (x => 440, y => 42),
  (x => 432, y => 43),
  (x => 433, y => 43),
  (x => 434, y => 43),
  (x => 435, y => 43),
  (x => 436, y => 43),
  (x => 437, y => 43),
  (x => 438, y => 43),
  (x => 439, y => 43),
  (x => 434, y => 44),
  (x => 435, y => 44),
  (x => 436, y => 44),
  (x => 437, y => 44)
);
constant p2_9: CoordPairArray(0 to 185) := (
  (x => 432, y => 22),
  (x => 433, y => 22),
  (x => 434, y => 22),
  (x => 435, y => 22),
  (x => 436, y => 22),
  (x => 437, y => 22),
  (x => 431, y => 23),
  (x => 432, y => 23),
  (x => 433, y => 23),
  (x => 434, y => 23),
  (x => 435, y => 23),
  (x => 436, y => 23),
  (x => 437, y => 23),
  (x => 438, y => 23),
  (x => 430, y => 24),
  (x => 431, y => 24),
  (x => 432, y => 24),
  (x => 433, y => 24),
  (x => 434, y => 24),
  (x => 435, y => 24),
  (x => 436, y => 24),
  (x => 437, y => 24),
  (x => 438, y => 24),
  (x => 439, y => 24),
  (x => 430, y => 25),
  (x => 431, y => 25),
  (x => 432, y => 25),
  (x => 433, y => 25),
  (x => 434, y => 25),
  (x => 435, y => 25),
  (x => 436, y => 25),
  (x => 437, y => 25),
  (x => 438, y => 25),
  (x => 439, y => 25),
  (x => 440, y => 25),
  (x => 430, y => 26),
  (x => 431, y => 26),
  (x => 432, y => 26),
  (x => 433, y => 26),
  (x => 437, y => 26),
  (x => 438, y => 26),
  (x => 439, y => 26),
  (x => 440, y => 26),
  (x => 429, y => 27),
  (x => 430, y => 27),
  (x => 431, y => 27),
  (x => 432, y => 27),
  (x => 437, y => 27),
  (x => 438, y => 27),
  (x => 439, y => 27),
  (x => 440, y => 27),
  (x => 429, y => 28),
  (x => 430, y => 28),
  (x => 431, y => 28),
  (x => 432, y => 28),
  (x => 438, y => 28),
  (x => 439, y => 28),
  (x => 440, y => 28),
  (x => 429, y => 29),
  (x => 430, y => 29),
  (x => 431, y => 29),
  (x => 432, y => 29),
  (x => 438, y => 29),
  (x => 439, y => 29),
  (x => 440, y => 29),
  (x => 441, y => 29),
  (x => 429, y => 30),
  (x => 430, y => 30),
  (x => 431, y => 30),
  (x => 432, y => 30),
  (x => 438, y => 30),
  (x => 439, y => 30),
  (x => 440, y => 30),
  (x => 441, y => 30),
  (x => 429, y => 31),
  (x => 430, y => 31),
  (x => 431, y => 31),
  (x => 432, y => 31),
  (x => 437, y => 31),
  (x => 438, y => 31),
  (x => 439, y => 31),
  (x => 440, y => 31),
  (x => 441, y => 31),
  (x => 429, y => 32),
  (x => 430, y => 32),
  (x => 431, y => 32),
  (x => 432, y => 32),
  (x => 433, y => 32),
  (x => 437, y => 32),
  (x => 438, y => 32),
  (x => 439, y => 32),
  (x => 440, y => 32),
  (x => 441, y => 32),
  (x => 430, y => 33),
  (x => 431, y => 33),
  (x => 432, y => 33),
  (x => 433, y => 33),
  (x => 434, y => 33),
  (x => 435, y => 33),
  (x => 436, y => 33),
  (x => 437, y => 33),
  (x => 438, y => 33),
  (x => 439, y => 33),
  (x => 440, y => 33),
  (x => 441, y => 33),
  (x => 430, y => 34),
  (x => 431, y => 34),
  (x => 432, y => 34),
  (x => 433, y => 34),
  (x => 434, y => 34),
  (x => 435, y => 34),
  (x => 436, y => 34),
  (x => 437, y => 34),
  (x => 438, y => 34),
  (x => 439, y => 34),
  (x => 440, y => 34),
  (x => 441, y => 34),
  (x => 431, y => 35),
  (x => 432, y => 35),
  (x => 433, y => 35),
  (x => 434, y => 35),
  (x => 435, y => 35),
  (x => 438, y => 35),
  (x => 439, y => 35),
  (x => 440, y => 35),
  (x => 441, y => 35),
  (x => 433, y => 36),
  (x => 434, y => 36),
  (x => 438, y => 36),
  (x => 439, y => 36),
  (x => 440, y => 36),
  (x => 441, y => 36),
  (x => 438, y => 37),
  (x => 439, y => 37),
  (x => 440, y => 37),
  (x => 441, y => 37),
  (x => 438, y => 38),
  (x => 439, y => 38),
  (x => 440, y => 38),
  (x => 437, y => 39),
  (x => 438, y => 39),
  (x => 439, y => 39),
  (x => 440, y => 39),
  (x => 437, y => 40),
  (x => 438, y => 40),
  (x => 439, y => 40),
  (x => 440, y => 40),
  (x => 435, y => 41),
  (x => 436, y => 41),
  (x => 437, y => 41),
  (x => 438, y => 41),
  (x => 439, y => 41),
  (x => 430, y => 42),
  (x => 431, y => 42),
  (x => 432, y => 42),
  (x => 433, y => 42),
  (x => 434, y => 42),
  (x => 435, y => 42),
  (x => 436, y => 42),
  (x => 437, y => 42),
  (x => 438, y => 42),
  (x => 439, y => 42),
  (x => 430, y => 43),
  (x => 431, y => 43),
  (x => 432, y => 43),
  (x => 433, y => 43),
  (x => 434, y => 43),
  (x => 435, y => 43),
  (x => 436, y => 43),
  (x => 437, y => 43),
  (x => 438, y => 43),
  (x => 430, y => 44),
  (x => 431, y => 44),
  (x => 432, y => 44),
  (x => 433, y => 44),
  (x => 434, y => 44),
  (x => 435, y => 44),
  (x => 436, y => 44),
  (x => 437, y => 44),
  (x => 430, y => 45),
  (x => 431, y => 45),
  (x => 432, y => 45),
  (x => 433, y => 45),
  (x => 434, y => 45),
  (x => 435, y => 45),
  (x => 436, y => 45)
);
	
	
end TXT_LIB;